module InvAES_S(
  input        clock,
  input        reset,
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _GEN_1 = 4'h0 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h9 : 8'h52; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_2 = 4'h0 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h6a : _GEN_1; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_3 = 4'h0 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hd5 : _GEN_2; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_4 = 4'h0 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h30 : _GEN_3; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_5 = 4'h0 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h36 : _GEN_4; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_6 = 4'h0 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'ha5 : _GEN_5; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_7 = 4'h0 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h38 : _GEN_6; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_8 = 4'h0 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hbf : _GEN_7; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_9 = 4'h0 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h40 : _GEN_8; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_10 = 4'h0 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'ha3 : _GEN_9; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_11 = 4'h0 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h9e : _GEN_10; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_12 = 4'h0 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h81 : _GEN_11; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_13 = 4'h0 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hf3 : _GEN_12; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_14 = 4'h0 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hd7 : _GEN_13; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_15 = 4'h0 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hfb : _GEN_14; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_16 = 4'h1 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h7c : _GEN_15; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_17 = 4'h1 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'he3 : _GEN_16; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_18 = 4'h1 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h39 : _GEN_17; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_19 = 4'h1 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h82 : _GEN_18; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_20 = 4'h1 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h9b : _GEN_19; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_21 = 4'h1 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h2f : _GEN_20; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_22 = 4'h1 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hff : _GEN_21; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_23 = 4'h1 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h87 : _GEN_22; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_24 = 4'h1 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h34 : _GEN_23; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_25 = 4'h1 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h8e : _GEN_24; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_26 = 4'h1 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h43 : _GEN_25; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_27 = 4'h1 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h44 : _GEN_26; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_28 = 4'h1 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hc4 : _GEN_27; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_29 = 4'h1 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hde : _GEN_28; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_30 = 4'h1 == io_in[7:4] & 4'he == io_in[3:0] ? 8'he9 : _GEN_29; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_31 = 4'h1 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hcb : _GEN_30; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_32 = 4'h2 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h54 : _GEN_31; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_33 = 4'h2 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h7b : _GEN_32; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_34 = 4'h2 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h94 : _GEN_33; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_35 = 4'h2 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h32 : _GEN_34; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_36 = 4'h2 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'ha6 : _GEN_35; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_37 = 4'h2 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hc2 : _GEN_36; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_38 = 4'h2 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h23 : _GEN_37; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_39 = 4'h2 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h3d : _GEN_38; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_40 = 4'h2 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hee : _GEN_39; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_41 = 4'h2 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h4c : _GEN_40; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_42 = 4'h2 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h95 : _GEN_41; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_43 = 4'h2 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hb : _GEN_42; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_44 = 4'h2 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h42 : _GEN_43; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_45 = 4'h2 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hfa : _GEN_44; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_46 = 4'h2 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hc3 : _GEN_45; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_47 = 4'h2 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h4e : _GEN_46; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_48 = 4'h3 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h8 : _GEN_47; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_49 = 4'h3 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h2e : _GEN_48; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_50 = 4'h3 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'ha1 : _GEN_49; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_51 = 4'h3 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h66 : _GEN_50; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_52 = 4'h3 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h28 : _GEN_51; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_53 = 4'h3 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hd9 : _GEN_52; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_54 = 4'h3 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h24 : _GEN_53; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_55 = 4'h3 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hb2 : _GEN_54; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_56 = 4'h3 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h76 : _GEN_55; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_57 = 4'h3 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h5b : _GEN_56; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_58 = 4'h3 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'ha2 : _GEN_57; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_59 = 4'h3 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h49 : _GEN_58; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_60 = 4'h3 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h6d : _GEN_59; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_61 = 4'h3 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h8b : _GEN_60; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_62 = 4'h3 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hd1 : _GEN_61; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_63 = 4'h3 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h25 : _GEN_62; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_64 = 4'h4 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h72 : _GEN_63; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_65 = 4'h4 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hf8 : _GEN_64; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_66 = 4'h4 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'hf6 : _GEN_65; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_67 = 4'h4 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h64 : _GEN_66; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_68 = 4'h4 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h86 : _GEN_67; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_69 = 4'h4 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h68 : _GEN_68; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_70 = 4'h4 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h98 : _GEN_69; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_71 = 4'h4 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h16 : _GEN_70; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_72 = 4'h4 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hd4 : _GEN_71; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_73 = 4'h4 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'ha4 : _GEN_72; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_74 = 4'h4 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h5c : _GEN_73; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_75 = 4'h4 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hcc : _GEN_74; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_76 = 4'h4 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h5d : _GEN_75; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_77 = 4'h4 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h65 : _GEN_76; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_78 = 4'h4 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hb6 : _GEN_77; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_79 = 4'h4 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h92 : _GEN_78; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_80 = 4'h5 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h6c : _GEN_79; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_81 = 4'h5 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h70 : _GEN_80; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_82 = 4'h5 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h48 : _GEN_81; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_83 = 4'h5 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h50 : _GEN_82; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_84 = 4'h5 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hfd : _GEN_83; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_85 = 4'h5 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hed : _GEN_84; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_86 = 4'h5 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hb9 : _GEN_85; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_87 = 4'h5 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hda : _GEN_86; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_88 = 4'h5 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h5e : _GEN_87; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_89 = 4'h5 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h15 : _GEN_88; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_90 = 4'h5 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h46 : _GEN_89; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_91 = 4'h5 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h57 : _GEN_90; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_92 = 4'h5 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'ha7 : _GEN_91; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_93 = 4'h5 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h8d : _GEN_92; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_94 = 4'h5 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h9d : _GEN_93; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_95 = 4'h5 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h84 : _GEN_94; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_96 = 4'h6 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h90 : _GEN_95; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_97 = 4'h6 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hd8 : _GEN_96; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_98 = 4'h6 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'hab : _GEN_97; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_99 = 4'h6 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h0 : _GEN_98; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_100 = 4'h6 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h8c : _GEN_99; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_101 = 4'h6 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hbc : _GEN_100; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_102 = 4'h6 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hd3 : _GEN_101; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_103 = 4'h6 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'ha : _GEN_102; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_104 = 4'h6 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hf7 : _GEN_103; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_105 = 4'h6 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'he4 : _GEN_104; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_106 = 4'h6 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h58 : _GEN_105; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_107 = 4'h6 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h5 : _GEN_106; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_108 = 4'h6 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hb8 : _GEN_107; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_109 = 4'h6 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hb3 : _GEN_108; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_110 = 4'h6 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h45 : _GEN_109; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_111 = 4'h6 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h6 : _GEN_110; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_112 = 4'h7 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hd0 : _GEN_111; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_113 = 4'h7 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h2c : _GEN_112; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_114 = 4'h7 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h1e : _GEN_113; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_115 = 4'h7 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h8f : _GEN_114; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_116 = 4'h7 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hca : _GEN_115; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_117 = 4'h7 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h3f : _GEN_116; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_118 = 4'h7 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hf : _GEN_117; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_119 = 4'h7 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h2 : _GEN_118; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_120 = 4'h7 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hc1 : _GEN_119; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_121 = 4'h7 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'haf : _GEN_120; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_122 = 4'h7 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hbd : _GEN_121; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_123 = 4'h7 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h3 : _GEN_122; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_124 = 4'h7 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h1 : _GEN_123; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_125 = 4'h7 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h13 : _GEN_124; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_126 = 4'h7 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h8a : _GEN_125; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_127 = 4'h7 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h6b : _GEN_126; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_128 = 4'h8 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h3a : _GEN_127; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_129 = 4'h8 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h91 : _GEN_128; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_130 = 4'h8 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h11 : _GEN_129; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_131 = 4'h8 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h41 : _GEN_130; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_132 = 4'h8 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h4f : _GEN_131; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_133 = 4'h8 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h67 : _GEN_132; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_134 = 4'h8 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hdc : _GEN_133; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_135 = 4'h8 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hea : _GEN_134; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_136 = 4'h8 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h97 : _GEN_135; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_137 = 4'h8 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hf2 : _GEN_136; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_138 = 4'h8 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hcf : _GEN_137; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_139 = 4'h8 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hce : _GEN_138; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_140 = 4'h8 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hf0 : _GEN_139; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_141 = 4'h8 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hb4 : _GEN_140; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_142 = 4'h8 == io_in[7:4] & 4'he == io_in[3:0] ? 8'he6 : _GEN_141; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_143 = 4'h8 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h73 : _GEN_142; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_144 = 4'h9 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h96 : _GEN_143; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_145 = 4'h9 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hac : _GEN_144; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_146 = 4'h9 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h74 : _GEN_145; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_147 = 4'h9 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h22 : _GEN_146; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_148 = 4'h9 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'he7 : _GEN_147; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_149 = 4'h9 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'had : _GEN_148; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_150 = 4'h9 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h35 : _GEN_149; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_151 = 4'h9 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h85 : _GEN_150; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_152 = 4'h9 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'he2 : _GEN_151; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_153 = 4'h9 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hf9 : _GEN_152; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_154 = 4'h9 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h37 : _GEN_153; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_155 = 4'h9 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'he8 : _GEN_154; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_156 = 4'h9 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h1c : _GEN_155; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_157 = 4'h9 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h75 : _GEN_156; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_158 = 4'h9 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hdf : _GEN_157; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_159 = 4'h9 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h6e : _GEN_158; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_160 = 4'ha == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h47 : _GEN_159; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_161 = 4'ha == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hf1 : _GEN_160; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_162 = 4'ha == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h1a : _GEN_161; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_163 = 4'ha == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h71 : _GEN_162; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_164 = 4'ha == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h1d : _GEN_163; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_165 = 4'ha == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h29 : _GEN_164; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_166 = 4'ha == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hc5 : _GEN_165; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_167 = 4'ha == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h89 : _GEN_166; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_168 = 4'ha == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h6f : _GEN_167; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_169 = 4'ha == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hb7 : _GEN_168; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_170 = 4'ha == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h62 : _GEN_169; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_171 = 4'ha == io_in[7:4] & 4'hb == io_in[3:0] ? 8'he : _GEN_170; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_172 = 4'ha == io_in[7:4] & 4'hc == io_in[3:0] ? 8'haa : _GEN_171; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_173 = 4'ha == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h18 : _GEN_172; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_174 = 4'ha == io_in[7:4] & 4'he == io_in[3:0] ? 8'hbe : _GEN_173; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_175 = 4'ha == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h1b : _GEN_174; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_176 = 4'hb == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hfc : _GEN_175; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_177 = 4'hb == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h56 : _GEN_176; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_178 = 4'hb == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h3e : _GEN_177; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_179 = 4'hb == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h4b : _GEN_178; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_180 = 4'hb == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hc6 : _GEN_179; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_181 = 4'hb == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hd2 : _GEN_180; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_182 = 4'hb == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h79 : _GEN_181; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_183 = 4'hb == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h20 : _GEN_182; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_184 = 4'hb == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h9a : _GEN_183; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_185 = 4'hb == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hdb : _GEN_184; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_186 = 4'hb == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hc0 : _GEN_185; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_187 = 4'hb == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hfe : _GEN_186; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_188 = 4'hb == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h78 : _GEN_187; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_189 = 4'hb == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hcd : _GEN_188; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_190 = 4'hb == io_in[7:4] & 4'he == io_in[3:0] ? 8'h5a : _GEN_189; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_191 = 4'hb == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hf4 : _GEN_190; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_192 = 4'hc == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h1f : _GEN_191; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_193 = 4'hc == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hdd : _GEN_192; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_194 = 4'hc == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'ha8 : _GEN_193; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_195 = 4'hc == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h33 : _GEN_194; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_196 = 4'hc == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h88 : _GEN_195; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_197 = 4'hc == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h7 : _GEN_196; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_198 = 4'hc == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hc7 : _GEN_197; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_199 = 4'hc == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h31 : _GEN_198; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_200 = 4'hc == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hb1 : _GEN_199; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_201 = 4'hc == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h12 : _GEN_200; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_202 = 4'hc == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h10 : _GEN_201; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_203 = 4'hc == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h59 : _GEN_202; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_204 = 4'hc == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h27 : _GEN_203; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_205 = 4'hc == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h80 : _GEN_204; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_206 = 4'hc == io_in[7:4] & 4'he == io_in[3:0] ? 8'hec : _GEN_205; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_207 = 4'hc == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h5f : _GEN_206; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_208 = 4'hd == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h60 : _GEN_207; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_209 = 4'hd == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h51 : _GEN_208; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_210 = 4'hd == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h7f : _GEN_209; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_211 = 4'hd == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'ha9 : _GEN_210; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_212 = 4'hd == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h19 : _GEN_211; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_213 = 4'hd == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hb5 : _GEN_212; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_214 = 4'hd == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h4a : _GEN_213; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_215 = 4'hd == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hd : _GEN_214; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_216 = 4'hd == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h2d : _GEN_215; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_217 = 4'hd == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'he5 : _GEN_216; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_218 = 4'hd == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h7a : _GEN_217; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_219 = 4'hd == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h9f : _GEN_218; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_220 = 4'hd == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h93 : _GEN_219; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_221 = 4'hd == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hc9 : _GEN_220; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_222 = 4'hd == io_in[7:4] & 4'he == io_in[3:0] ? 8'h9c : _GEN_221; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_223 = 4'hd == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hef : _GEN_222; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_224 = 4'he == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'ha0 : _GEN_223; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_225 = 4'he == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'he0 : _GEN_224; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_226 = 4'he == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h3b : _GEN_225; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_227 = 4'he == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h4d : _GEN_226; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_228 = 4'he == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hae : _GEN_227; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_229 = 4'he == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h2a : _GEN_228; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_230 = 4'he == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hf5 : _GEN_229; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_231 = 4'he == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hb0 : _GEN_230; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_232 = 4'he == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hc8 : _GEN_231; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_233 = 4'he == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'heb : _GEN_232; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_234 = 4'he == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hbb : _GEN_233; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_235 = 4'he == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h3c : _GEN_234; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_236 = 4'he == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h83 : _GEN_235; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_237 = 4'he == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h53 : _GEN_236; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_238 = 4'he == io_in[7:4] & 4'he == io_in[3:0] ? 8'h99 : _GEN_237; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_239 = 4'he == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h61 : _GEN_238; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_240 = 4'hf == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h17 : _GEN_239; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_241 = 4'hf == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h2b : _GEN_240; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_242 = 4'hf == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h4 : _GEN_241; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_243 = 4'hf == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h7e : _GEN_242; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_244 = 4'hf == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hba : _GEN_243; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_245 = 4'hf == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h77 : _GEN_244; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_246 = 4'hf == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hd6 : _GEN_245; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_247 = 4'hf == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h26 : _GEN_246; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_248 = 4'hf == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'he1 : _GEN_247; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_249 = 4'hf == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h69 : _GEN_248; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_250 = 4'hf == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h14 : _GEN_249; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_251 = 4'hf == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h63 : _GEN_250; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_252 = 4'hf == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h55 : _GEN_251; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_253 = 4'hf == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h21 : _GEN_252; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  wire [7:0] _GEN_254 = 4'hf == io_in[7:4] & 4'he == io_in[3:0] ? 8'hc : _GEN_253; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
  assign io_out = 4'hf == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h7d : _GEN_254; // @[AES_Pipelined.scala 270:10 AES_Pipelined.scala 270:10]
endmodule
