module AES_InitialOperation(
  input  [127:0] io_text,
  input  [127:0] io_key,
  output [7:0]   io_out_state_0_0,
  output [7:0]   io_out_state_0_1,
  output [7:0]   io_out_state_0_2,
  output [7:0]   io_out_state_0_3,
  output [7:0]   io_out_state_1_0,
  output [7:0]   io_out_state_1_1,
  output [7:0]   io_out_state_1_2,
  output [7:0]   io_out_state_1_3,
  output [7:0]   io_out_state_2_0,
  output [7:0]   io_out_state_2_1,
  output [7:0]   io_out_state_2_2,
  output [7:0]   io_out_state_2_3,
  output [7:0]   io_out_state_3_0,
  output [7:0]   io_out_state_3_1,
  output [7:0]   io_out_state_3_2,
  output [7:0]   io_out_state_3_3,
  output [7:0]   io_out_key_0_0,
  output [7:0]   io_out_key_0_1,
  output [7:0]   io_out_key_0_2,
  output [7:0]   io_out_key_0_3,
  output [7:0]   io_out_key_1_0,
  output [7:0]   io_out_key_1_1,
  output [7:0]   io_out_key_1_2,
  output [7:0]   io_out_key_1_3,
  output [7:0]   io_out_key_2_0,
  output [7:0]   io_out_key_2_1,
  output [7:0]   io_out_key_2_2,
  output [7:0]   io_out_key_2_3,
  output [7:0]   io_out_key_3_0,
  output [7:0]   io_out_key_3_1,
  output [7:0]   io_out_key_3_2,
  output [7:0]   io_out_key_3_3
);
  assign io_out_state_0_0 = io_text[127:120]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_0_1 = io_text[119:112]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_0_2 = io_text[111:104]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_0_3 = io_text[103:96]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_1_0 = io_text[95:88]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_1_1 = io_text[87:80]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_1_2 = io_text[79:72]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_1_3 = io_text[71:64]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_2_0 = io_text[63:56]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_2_1 = io_text[55:48]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_2_2 = io_text[47:40]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_2_3 = io_text[39:32]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_3_0 = io_text[31:24]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_3_1 = io_text[23:16]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_3_2 = io_text[15:8]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_state_3_3 = io_text[7:0]; // @[AES_EncryptionFSM.scala 80:40]
  assign io_out_key_0_0 = io_key[127:120]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_0_1 = io_key[119:112]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_0_2 = io_key[111:104]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_0_3 = io_key[103:96]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_1_0 = io_key[95:88]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_1_1 = io_key[87:80]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_1_2 = io_key[79:72]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_1_3 = io_key[71:64]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_2_0 = io_key[63:56]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_2_1 = io_key[55:48]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_2_2 = io_key[47:40]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_2_3 = io_key[39:32]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_3_0 = io_key[31:24]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_3_1 = io_key[23:16]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_3_2 = io_key[15:8]; // @[AES_EncryptionFSM.scala 81:37]
  assign io_out_key_3_3 = io_key[7:0]; // @[AES_EncryptionFSM.scala 81:37]
endmodule
module AES_FinalOperation(
  output [127:0] io_out_text,
  output [127:0] io_out_key,
  input  [7:0]   io_in_state_0_0,
  input  [7:0]   io_in_state_0_1,
  input  [7:0]   io_in_state_0_2,
  input  [7:0]   io_in_state_0_3,
  input  [7:0]   io_in_state_1_0,
  input  [7:0]   io_in_state_1_1,
  input  [7:0]   io_in_state_1_2,
  input  [7:0]   io_in_state_1_3,
  input  [7:0]   io_in_state_2_0,
  input  [7:0]   io_in_state_2_1,
  input  [7:0]   io_in_state_2_2,
  input  [7:0]   io_in_state_2_3,
  input  [7:0]   io_in_state_3_0,
  input  [7:0]   io_in_state_3_1,
  input  [7:0]   io_in_state_3_2,
  input  [7:0]   io_in_state_3_3,
  input  [7:0]   io_in_key_0_0,
  input  [7:0]   io_in_key_0_1,
  input  [7:0]   io_in_key_0_2,
  input  [7:0]   io_in_key_0_3,
  input  [7:0]   io_in_key_1_0,
  input  [7:0]   io_in_key_1_1,
  input  [7:0]   io_in_key_1_2,
  input  [7:0]   io_in_key_1_3,
  input  [7:0]   io_in_key_2_0,
  input  [7:0]   io_in_key_2_1,
  input  [7:0]   io_in_key_2_2,
  input  [7:0]   io_in_key_2_3,
  input  [7:0]   io_in_key_3_0,
  input  [7:0]   io_in_key_3_1,
  input  [7:0]   io_in_key_3_2,
  input  [7:0]   io_in_key_3_3
);
  wire [7:0] hi_hi_hi_hi = io_in_state_0_0 ^ io_in_key_0_0; // @[AES_EncryptionFSM.scala 93:39]
  wire [7:0] hi_hi_hi_lo = io_in_state_0_1 ^ io_in_key_0_1; // @[AES_EncryptionFSM.scala 93:73]
  wire [7:0] hi_hi_lo_hi = io_in_state_0_2 ^ io_in_key_0_2; // @[AES_EncryptionFSM.scala 94:22]
  wire [7:0] hi_hi_lo_lo = io_in_state_0_3 ^ io_in_key_0_3; // @[AES_EncryptionFSM.scala 94:56]
  wire [7:0] hi_lo_hi_hi = io_in_state_1_0 ^ io_in_key_1_0; // @[AES_EncryptionFSM.scala 95:22]
  wire [7:0] hi_lo_hi_lo = io_in_state_1_1 ^ io_in_key_1_1; // @[AES_EncryptionFSM.scala 95:56]
  wire [7:0] hi_lo_lo_hi = io_in_state_1_2 ^ io_in_key_1_2; // @[AES_EncryptionFSM.scala 96:22]
  wire [7:0] hi_lo_lo_lo = io_in_state_1_3 ^ io_in_key_1_3; // @[AES_EncryptionFSM.scala 96:56]
  wire [7:0] lo_hi_hi_hi = io_in_state_2_0 ^ io_in_key_2_0; // @[AES_EncryptionFSM.scala 97:22]
  wire [7:0] lo_hi_hi_lo = io_in_state_2_1 ^ io_in_key_2_1; // @[AES_EncryptionFSM.scala 97:56]
  wire [7:0] lo_hi_lo_hi = io_in_state_2_2 ^ io_in_key_2_2; // @[AES_EncryptionFSM.scala 98:22]
  wire [7:0] lo_hi_lo_lo = io_in_state_2_3 ^ io_in_key_2_3; // @[AES_EncryptionFSM.scala 98:56]
  wire [7:0] lo_lo_hi_hi = io_in_state_3_0 ^ io_in_key_3_0; // @[AES_EncryptionFSM.scala 99:22]
  wire [7:0] lo_lo_hi_lo = io_in_state_3_1 ^ io_in_key_3_1; // @[AES_EncryptionFSM.scala 99:56]
  wire [7:0] lo_lo_lo_hi = io_in_state_3_2 ^ io_in_key_3_2; // @[AES_EncryptionFSM.scala 100:22]
  wire [7:0] lo_lo_lo_lo = io_in_state_3_3 ^ io_in_key_3_3; // @[AES_EncryptionFSM.scala 100:56]
  wire [63:0] lo = {lo_hi_hi_hi,lo_hi_hi_lo,lo_hi_lo_hi,lo_hi_lo_lo,lo_lo_hi_hi,lo_lo_hi_lo,lo_lo_lo_hi,lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] hi = {hi_hi_hi_hi,hi_hi_hi_lo,hi_hi_lo_hi,hi_hi_lo_lo,hi_lo_hi_hi,hi_lo_hi_lo,hi_lo_lo_hi,hi_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] lo_1 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3,io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,
    io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [63:0] hi_1 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3,io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,
    io_in_key_1_3}; // @[Cat.scala 30:58]
  assign io_out_text = {hi,lo}; // @[Cat.scala 30:58]
  assign io_out_key = {hi_1,lo_1}; // @[Cat.scala 30:58]
endmodule
module AES_S(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _GEN_1 = 4'h0 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h7c : 8'h63; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_2 = 4'h0 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h77 : _GEN_1; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_3 = 4'h0 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h7b : _GEN_2; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_4 = 4'h0 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hf2 : _GEN_3; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_5 = 4'h0 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h6b : _GEN_4; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_6 = 4'h0 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h6f : _GEN_5; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_7 = 4'h0 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hc5 : _GEN_6; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_8 = 4'h0 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h30 : _GEN_7; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_9 = 4'h0 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h1 : _GEN_8; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_10 = 4'h0 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h67 : _GEN_9; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_11 = 4'h0 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h2b : _GEN_10; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_12 = 4'h0 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hfe : _GEN_11; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_13 = 4'h0 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hd7 : _GEN_12; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_14 = 4'h0 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hab : _GEN_13; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_15 = 4'h0 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h76 : _GEN_14; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_16 = 4'h1 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hca : _GEN_15; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_17 = 4'h1 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h82 : _GEN_16; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_18 = 4'h1 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'hc9 : _GEN_17; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_19 = 4'h1 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h7d : _GEN_18; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_20 = 4'h1 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hfa : _GEN_19; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_21 = 4'h1 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h59 : _GEN_20; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_22 = 4'h1 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h47 : _GEN_21; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_23 = 4'h1 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hf0 : _GEN_22; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_24 = 4'h1 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'had : _GEN_23; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_25 = 4'h1 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hd4 : _GEN_24; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_26 = 4'h1 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'ha2 : _GEN_25; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_27 = 4'h1 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'haf : _GEN_26; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_28 = 4'h1 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h9c : _GEN_27; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_29 = 4'h1 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'ha4 : _GEN_28; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_30 = 4'h1 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h72 : _GEN_29; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_31 = 4'h1 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hc0 : _GEN_30; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_32 = 4'h2 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hb7 : _GEN_31; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_33 = 4'h2 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hfd : _GEN_32; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_34 = 4'h2 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h93 : _GEN_33; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_35 = 4'h2 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h26 : _GEN_34; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_36 = 4'h2 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h36 : _GEN_35; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_37 = 4'h2 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h3f : _GEN_36; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_38 = 4'h2 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hf7 : _GEN_37; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_39 = 4'h2 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hcc : _GEN_38; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_40 = 4'h2 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h34 : _GEN_39; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_41 = 4'h2 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'ha5 : _GEN_40; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_42 = 4'h2 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'he5 : _GEN_41; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_43 = 4'h2 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hf1 : _GEN_42; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_44 = 4'h2 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h71 : _GEN_43; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_45 = 4'h2 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hd8 : _GEN_44; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_46 = 4'h2 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h31 : _GEN_45; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_47 = 4'h2 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h15 : _GEN_46; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_48 = 4'h3 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h4 : _GEN_47; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_49 = 4'h3 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hc7 : _GEN_48; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_50 = 4'h3 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h23 : _GEN_49; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_51 = 4'h3 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hc3 : _GEN_50; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_52 = 4'h3 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h18 : _GEN_51; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_53 = 4'h3 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h96 : _GEN_52; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_54 = 4'h3 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h5 : _GEN_53; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_55 = 4'h3 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h9a : _GEN_54; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_56 = 4'h3 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h7 : _GEN_55; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_57 = 4'h3 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h12 : _GEN_56; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_58 = 4'h3 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h80 : _GEN_57; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_59 = 4'h3 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'he2 : _GEN_58; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_60 = 4'h3 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'heb : _GEN_59; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_61 = 4'h3 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h27 : _GEN_60; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_62 = 4'h3 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hb2 : _GEN_61; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_63 = 4'h3 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h75 : _GEN_62; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_64 = 4'h4 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h9 : _GEN_63; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_65 = 4'h4 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h83 : _GEN_64; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_66 = 4'h4 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h2c : _GEN_65; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_67 = 4'h4 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h1a : _GEN_66; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_68 = 4'h4 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h1b : _GEN_67; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_69 = 4'h4 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h6e : _GEN_68; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_70 = 4'h4 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h5a : _GEN_69; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_71 = 4'h4 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'ha0 : _GEN_70; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_72 = 4'h4 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h52 : _GEN_71; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_73 = 4'h4 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h3b : _GEN_72; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_74 = 4'h4 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hd6 : _GEN_73; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_75 = 4'h4 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hb3 : _GEN_74; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_76 = 4'h4 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h29 : _GEN_75; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_77 = 4'h4 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'he3 : _GEN_76; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_78 = 4'h4 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h2f : _GEN_77; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_79 = 4'h4 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h84 : _GEN_78; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_80 = 4'h5 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h53 : _GEN_79; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_81 = 4'h5 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hd1 : _GEN_80; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_82 = 4'h5 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h0 : _GEN_81; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_83 = 4'h5 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hed : _GEN_82; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_84 = 4'h5 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h20 : _GEN_83; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_85 = 4'h5 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hfc : _GEN_84; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_86 = 4'h5 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hb1 : _GEN_85; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_87 = 4'h5 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h5b : _GEN_86; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_88 = 4'h5 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h6a : _GEN_87; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_89 = 4'h5 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hcb : _GEN_88; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_90 = 4'h5 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hbe : _GEN_89; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_91 = 4'h5 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h39 : _GEN_90; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_92 = 4'h5 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h4a : _GEN_91; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_93 = 4'h5 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h4c : _GEN_92; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_94 = 4'h5 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h58 : _GEN_93; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_95 = 4'h5 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hcf : _GEN_94; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_96 = 4'h6 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hd0 : _GEN_95; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_97 = 4'h6 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hef : _GEN_96; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_98 = 4'h6 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'haa : _GEN_97; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_99 = 4'h6 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hfb : _GEN_98; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_100 = 4'h6 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h43 : _GEN_99; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_101 = 4'h6 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h4d : _GEN_100; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_102 = 4'h6 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h33 : _GEN_101; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_103 = 4'h6 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h85 : _GEN_102; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_104 = 4'h6 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h45 : _GEN_103; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_105 = 4'h6 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hf9 : _GEN_104; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_106 = 4'h6 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h2 : _GEN_105; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_107 = 4'h6 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h7f : _GEN_106; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_108 = 4'h6 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h50 : _GEN_107; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_109 = 4'h6 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h3c : _GEN_108; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_110 = 4'h6 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h9f : _GEN_109; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_111 = 4'h6 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'ha8 : _GEN_110; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_112 = 4'h7 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h51 : _GEN_111; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_113 = 4'h7 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'ha3 : _GEN_112; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_114 = 4'h7 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h40 : _GEN_113; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_115 = 4'h7 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h8f : _GEN_114; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_116 = 4'h7 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h92 : _GEN_115; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_117 = 4'h7 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h9d : _GEN_116; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_118 = 4'h7 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h38 : _GEN_117; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_119 = 4'h7 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hf5 : _GEN_118; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_120 = 4'h7 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hbc : _GEN_119; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_121 = 4'h7 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hb6 : _GEN_120; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_122 = 4'h7 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hda : _GEN_121; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_123 = 4'h7 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h21 : _GEN_122; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_124 = 4'h7 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h10 : _GEN_123; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_125 = 4'h7 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hff : _GEN_124; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_126 = 4'h7 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hf3 : _GEN_125; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_127 = 4'h7 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hd2 : _GEN_126; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_128 = 4'h8 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hcd : _GEN_127; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_129 = 4'h8 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hc : _GEN_128; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_130 = 4'h8 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h13 : _GEN_129; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_131 = 4'h8 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hec : _GEN_130; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_132 = 4'h8 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h5f : _GEN_131; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_133 = 4'h8 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h97 : _GEN_132; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_134 = 4'h8 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h44 : _GEN_133; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_135 = 4'h8 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h17 : _GEN_134; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_136 = 4'h8 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hc4 : _GEN_135; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_137 = 4'h8 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'ha7 : _GEN_136; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_138 = 4'h8 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h7e : _GEN_137; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_139 = 4'h8 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h3d : _GEN_138; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_140 = 4'h8 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h64 : _GEN_139; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_141 = 4'h8 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h5d : _GEN_140; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_142 = 4'h8 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h19 : _GEN_141; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_143 = 4'h8 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h73 : _GEN_142; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_144 = 4'h9 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h60 : _GEN_143; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_145 = 4'h9 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h81 : _GEN_144; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_146 = 4'h9 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h4f : _GEN_145; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_147 = 4'h9 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hdc : _GEN_146; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_148 = 4'h9 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h22 : _GEN_147; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_149 = 4'h9 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h2a : _GEN_148; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_150 = 4'h9 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h90 : _GEN_149; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_151 = 4'h9 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h88 : _GEN_150; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_152 = 4'h9 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h46 : _GEN_151; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_153 = 4'h9 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hee : _GEN_152; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_154 = 4'h9 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hb8 : _GEN_153; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_155 = 4'h9 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h14 : _GEN_154; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_156 = 4'h9 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hde : _GEN_155; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_157 = 4'h9 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h5e : _GEN_156; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_158 = 4'h9 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hb : _GEN_157; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_159 = 4'h9 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hdb : _GEN_158; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_160 = 4'ha == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'he0 : _GEN_159; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_161 = 4'ha == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h32 : _GEN_160; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_162 = 4'ha == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h3a : _GEN_161; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_163 = 4'ha == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'ha : _GEN_162; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_164 = 4'ha == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h49 : _GEN_163; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_165 = 4'ha == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h6 : _GEN_164; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_166 = 4'ha == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h24 : _GEN_165; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_167 = 4'ha == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h5c : _GEN_166; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_168 = 4'ha == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hc2 : _GEN_167; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_169 = 4'ha == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hd3 : _GEN_168; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_170 = 4'ha == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hac : _GEN_169; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_171 = 4'ha == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h62 : _GEN_170; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_172 = 4'ha == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h91 : _GEN_171; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_173 = 4'ha == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h95 : _GEN_172; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_174 = 4'ha == io_in[7:4] & 4'he == io_in[3:0] ? 8'he4 : _GEN_173; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_175 = 4'ha == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h79 : _GEN_174; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_176 = 4'hb == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'he7 : _GEN_175; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_177 = 4'hb == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hc8 : _GEN_176; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_178 = 4'hb == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h37 : _GEN_177; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_179 = 4'hb == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h6d : _GEN_178; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_180 = 4'hb == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h8d : _GEN_179; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_181 = 4'hb == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hd5 : _GEN_180; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_182 = 4'hb == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h4e : _GEN_181; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_183 = 4'hb == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'ha9 : _GEN_182; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_184 = 4'hb == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h6c : _GEN_183; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_185 = 4'hb == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h56 : _GEN_184; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_186 = 4'hb == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hf4 : _GEN_185; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_187 = 4'hb == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hea : _GEN_186; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_188 = 4'hb == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h65 : _GEN_187; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_189 = 4'hb == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h7a : _GEN_188; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_190 = 4'hb == io_in[7:4] & 4'he == io_in[3:0] ? 8'hae : _GEN_189; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_191 = 4'hb == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h8 : _GEN_190; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_192 = 4'hc == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hba : _GEN_191; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_193 = 4'hc == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h78 : _GEN_192; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_194 = 4'hc == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h25 : _GEN_193; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_195 = 4'hc == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h2e : _GEN_194; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_196 = 4'hc == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h1c : _GEN_195; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_197 = 4'hc == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'ha6 : _GEN_196; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_198 = 4'hc == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hb4 : _GEN_197; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_199 = 4'hc == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hc6 : _GEN_198; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_200 = 4'hc == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'he8 : _GEN_199; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_201 = 4'hc == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hdd : _GEN_200; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_202 = 4'hc == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h74 : _GEN_201; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_203 = 4'hc == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h1f : _GEN_202; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_204 = 4'hc == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h4b : _GEN_203; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_205 = 4'hc == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hbd : _GEN_204; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_206 = 4'hc == io_in[7:4] & 4'he == io_in[3:0] ? 8'h8b : _GEN_205; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_207 = 4'hc == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h8a : _GEN_206; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_208 = 4'hd == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h70 : _GEN_207; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_209 = 4'hd == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h3e : _GEN_208; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_210 = 4'hd == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'hb5 : _GEN_209; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_211 = 4'hd == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h66 : _GEN_210; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_212 = 4'hd == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h48 : _GEN_211; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_213 = 4'hd == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h3 : _GEN_212; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_214 = 4'hd == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hf6 : _GEN_213; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_215 = 4'hd == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'he : _GEN_214; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_216 = 4'hd == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h61 : _GEN_215; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_217 = 4'hd == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h35 : _GEN_216; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_218 = 4'hd == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h57 : _GEN_217; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_219 = 4'hd == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hb9 : _GEN_218; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_220 = 4'hd == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h86 : _GEN_219; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_221 = 4'hd == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hc1 : _GEN_220; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_222 = 4'hd == io_in[7:4] & 4'he == io_in[3:0] ? 8'h1d : _GEN_221; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_223 = 4'hd == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h9e : _GEN_222; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_224 = 4'he == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'he1 : _GEN_223; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_225 = 4'he == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hf8 : _GEN_224; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_226 = 4'he == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h98 : _GEN_225; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_227 = 4'he == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h11 : _GEN_226; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_228 = 4'he == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h69 : _GEN_227; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_229 = 4'he == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hd9 : _GEN_228; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_230 = 4'he == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h8e : _GEN_229; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_231 = 4'he == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h94 : _GEN_230; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_232 = 4'he == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h9b : _GEN_231; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_233 = 4'he == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h1e : _GEN_232; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_234 = 4'he == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h87 : _GEN_233; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_235 = 4'he == io_in[7:4] & 4'hb == io_in[3:0] ? 8'he9 : _GEN_234; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_236 = 4'he == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hce : _GEN_235; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_237 = 4'he == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h55 : _GEN_236; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_238 = 4'he == io_in[7:4] & 4'he == io_in[3:0] ? 8'h28 : _GEN_237; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_239 = 4'he == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hdf : _GEN_238; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_240 = 4'hf == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h8c : _GEN_239; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_241 = 4'hf == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'ha1 : _GEN_240; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_242 = 4'hf == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h89 : _GEN_241; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_243 = 4'hf == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hd : _GEN_242; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_244 = 4'hf == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hbf : _GEN_243; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_245 = 4'hf == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'he6 : _GEN_244; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_246 = 4'hf == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h42 : _GEN_245; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_247 = 4'hf == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h68 : _GEN_246; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_248 = 4'hf == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h41 : _GEN_247; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_249 = 4'hf == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h99 : _GEN_248; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_250 = 4'hf == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h2d : _GEN_249; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_251 = 4'hf == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hf : _GEN_250; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_252 = 4'hf == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hb0 : _GEN_251; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_253 = 4'hf == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h54 : _GEN_252; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  wire [7:0] _GEN_254 = 4'hf == io_in[7:4] & 4'he == io_in[3:0] ? 8'hbb : _GEN_253; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
  assign io_out = 4'hf == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h16 : _GEN_254; // @[AES_EncryptionFSM.scala 394:10 AES_EncryptionFSM.scala 394:10]
endmodule
module AES_SubBytes(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3
);
  wire [7:0] PEs_0_0_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_0_0_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_0_1_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_0_1_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_0_2_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_0_2_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_0_3_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_0_3_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_1_0_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_1_0_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_1_1_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_1_1_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_1_2_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_1_2_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_1_3_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_1_3_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_2_0_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_2_0_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_2_1_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_2_1_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_2_2_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_2_2_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_2_3_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_2_3_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_3_0_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_3_0_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_3_1_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_3_1_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_3_2_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_3_2_io_out; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_3_3_io_in; // @[AES_EncryptionFSM.scala 341:22]
  wire [7:0] PEs_3_3_io_out; // @[AES_EncryptionFSM.scala 341:22]
  AES_S PEs_0_0 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_0_0_io_in),
    .io_out(PEs_0_0_io_out)
  );
  AES_S PEs_0_1 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_0_1_io_in),
    .io_out(PEs_0_1_io_out)
  );
  AES_S PEs_0_2 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_0_2_io_in),
    .io_out(PEs_0_2_io_out)
  );
  AES_S PEs_0_3 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_0_3_io_in),
    .io_out(PEs_0_3_io_out)
  );
  AES_S PEs_1_0 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_1_0_io_in),
    .io_out(PEs_1_0_io_out)
  );
  AES_S PEs_1_1 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_1_1_io_in),
    .io_out(PEs_1_1_io_out)
  );
  AES_S PEs_1_2 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_1_2_io_in),
    .io_out(PEs_1_2_io_out)
  );
  AES_S PEs_1_3 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_1_3_io_in),
    .io_out(PEs_1_3_io_out)
  );
  AES_S PEs_2_0 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_2_0_io_in),
    .io_out(PEs_2_0_io_out)
  );
  AES_S PEs_2_1 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_2_1_io_in),
    .io_out(PEs_2_1_io_out)
  );
  AES_S PEs_2_2 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_2_2_io_in),
    .io_out(PEs_2_2_io_out)
  );
  AES_S PEs_2_3 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_2_3_io_in),
    .io_out(PEs_2_3_io_out)
  );
  AES_S PEs_3_0 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_3_0_io_in),
    .io_out(PEs_3_0_io_out)
  );
  AES_S PEs_3_1 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_3_1_io_in),
    .io_out(PEs_3_1_io_out)
  );
  AES_S PEs_3_2 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_3_2_io_in),
    .io_out(PEs_3_2_io_out)
  );
  AES_S PEs_3_3 ( // @[AES_EncryptionFSM.scala 341:22]
    .io_in(PEs_3_3_io_in),
    .io_out(PEs_3_3_io_out)
  );
  assign io_out_state_0_0 = PEs_0_0_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_0_1 = PEs_0_1_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_0_2 = PEs_0_2_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_0_3 = PEs_0_3_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_1_0 = PEs_1_0_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_1_1 = PEs_1_1_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_1_2 = PEs_1_2_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_1_3 = PEs_1_3_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_2_0 = PEs_2_0_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_2_1 = PEs_2_1_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_2_2 = PEs_2_2_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_2_3 = PEs_2_3_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_3_0 = PEs_3_0_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_3_1 = PEs_3_1_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_3_2 = PEs_3_2_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign io_out_state_3_3 = PEs_3_3_io_out; // @[AES_EncryptionFSM.scala 350:26]
  assign PEs_0_0_io_in = io_in_state_0_0; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_0_1_io_in = io_in_state_0_1; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_0_2_io_in = io_in_state_0_2; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_0_3_io_in = io_in_state_0_3; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_1_0_io_in = io_in_state_1_0; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_1_1_io_in = io_in_state_1_1; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_1_2_io_in = io_in_state_1_2; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_1_3_io_in = io_in_state_1_3; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_2_0_io_in = io_in_state_2_0; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_2_1_io_in = io_in_state_2_1; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_2_2_io_in = io_in_state_2_2; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_2_3_io_in = io_in_state_2_3; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_3_0_io_in = io_in_state_3_0; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_3_1_io_in = io_in_state_3_1; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_3_2_io_in = io_in_state_3_2; // @[AES_EncryptionFSM.scala 349:23]
  assign PEs_3_3_io_in = io_in_state_3_3; // @[AES_EncryptionFSM.scala 349:23]
endmodule
module AES_ShiftRows(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3
);
  assign io_out_state_0_0 = io_in_state_0_0; // @[AES_EncryptionFSM.scala 310:22]
  assign io_out_state_0_1 = io_in_state_1_1; // @[AES_EncryptionFSM.scala 315:22]
  assign io_out_state_0_2 = io_in_state_2_2; // @[AES_EncryptionFSM.scala 320:22]
  assign io_out_state_0_3 = io_in_state_3_3; // @[AES_EncryptionFSM.scala 325:22]
  assign io_out_state_1_0 = io_in_state_1_0; // @[AES_EncryptionFSM.scala 311:22]
  assign io_out_state_1_1 = io_in_state_2_1; // @[AES_EncryptionFSM.scala 316:22]
  assign io_out_state_1_2 = io_in_state_3_2; // @[AES_EncryptionFSM.scala 321:22]
  assign io_out_state_1_3 = io_in_state_0_3; // @[AES_EncryptionFSM.scala 326:22]
  assign io_out_state_2_0 = io_in_state_2_0; // @[AES_EncryptionFSM.scala 312:22]
  assign io_out_state_2_1 = io_in_state_3_1; // @[AES_EncryptionFSM.scala 317:22]
  assign io_out_state_2_2 = io_in_state_0_2; // @[AES_EncryptionFSM.scala 322:22]
  assign io_out_state_2_3 = io_in_state_1_3; // @[AES_EncryptionFSM.scala 327:22]
  assign io_out_state_3_0 = io_in_state_3_0; // @[AES_EncryptionFSM.scala 313:22]
  assign io_out_state_3_1 = io_in_state_0_1; // @[AES_EncryptionFSM.scala 318:22]
  assign io_out_state_3_2 = io_in_state_1_2; // @[AES_EncryptionFSM.scala 323:22]
  assign io_out_state_3_3 = io_in_state_2_3; // @[AES_EncryptionFSM.scala 328:22]
endmodule
module AES_MixColumn(
  input  [7:0] io_in_0,
  input  [7:0] io_in_1,
  input  [7:0] io_in_2,
  input  [7:0] io_in_3,
  output [7:0] io_out_0,
  output [7:0] io_out_1,
  output [7:0] io_out_2,
  output [7:0] io_out_3
);
  wire [7:0] _GEN_1 = 8'h1 == io_in_0 ? 8'h2 : 8'h0; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_2 = 8'h2 == io_in_0 ? 8'h4 : _GEN_1; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_3 = 8'h3 == io_in_0 ? 8'h6 : _GEN_2; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_4 = 8'h4 == io_in_0 ? 8'h8 : _GEN_3; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_5 = 8'h5 == io_in_0 ? 8'ha : _GEN_4; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_6 = 8'h6 == io_in_0 ? 8'hc : _GEN_5; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_7 = 8'h7 == io_in_0 ? 8'he : _GEN_6; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_8 = 8'h8 == io_in_0 ? 8'h10 : _GEN_7; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_9 = 8'h9 == io_in_0 ? 8'h12 : _GEN_8; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_10 = 8'ha == io_in_0 ? 8'h14 : _GEN_9; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_11 = 8'hb == io_in_0 ? 8'h16 : _GEN_10; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_12 = 8'hc == io_in_0 ? 8'h18 : _GEN_11; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_13 = 8'hd == io_in_0 ? 8'h1a : _GEN_12; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_14 = 8'he == io_in_0 ? 8'h1c : _GEN_13; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_15 = 8'hf == io_in_0 ? 8'h1e : _GEN_14; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_16 = 8'h10 == io_in_0 ? 8'h20 : _GEN_15; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_17 = 8'h11 == io_in_0 ? 8'h22 : _GEN_16; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_18 = 8'h12 == io_in_0 ? 8'h24 : _GEN_17; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_19 = 8'h13 == io_in_0 ? 8'h26 : _GEN_18; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_20 = 8'h14 == io_in_0 ? 8'h28 : _GEN_19; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_21 = 8'h15 == io_in_0 ? 8'h2a : _GEN_20; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_22 = 8'h16 == io_in_0 ? 8'h2c : _GEN_21; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_23 = 8'h17 == io_in_0 ? 8'h2e : _GEN_22; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_24 = 8'h18 == io_in_0 ? 8'h30 : _GEN_23; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_25 = 8'h19 == io_in_0 ? 8'h32 : _GEN_24; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_26 = 8'h1a == io_in_0 ? 8'h34 : _GEN_25; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_27 = 8'h1b == io_in_0 ? 8'h36 : _GEN_26; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_28 = 8'h1c == io_in_0 ? 8'h38 : _GEN_27; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_29 = 8'h1d == io_in_0 ? 8'h3a : _GEN_28; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_30 = 8'h1e == io_in_0 ? 8'h3c : _GEN_29; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_31 = 8'h1f == io_in_0 ? 8'h3e : _GEN_30; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_32 = 8'h20 == io_in_0 ? 8'h40 : _GEN_31; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_33 = 8'h21 == io_in_0 ? 8'h42 : _GEN_32; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_34 = 8'h22 == io_in_0 ? 8'h44 : _GEN_33; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_35 = 8'h23 == io_in_0 ? 8'h46 : _GEN_34; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_36 = 8'h24 == io_in_0 ? 8'h48 : _GEN_35; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_37 = 8'h25 == io_in_0 ? 8'h4a : _GEN_36; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_38 = 8'h26 == io_in_0 ? 8'h4c : _GEN_37; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_39 = 8'h27 == io_in_0 ? 8'h4e : _GEN_38; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_40 = 8'h28 == io_in_0 ? 8'h50 : _GEN_39; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_41 = 8'h29 == io_in_0 ? 8'h52 : _GEN_40; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_42 = 8'h2a == io_in_0 ? 8'h54 : _GEN_41; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_43 = 8'h2b == io_in_0 ? 8'h56 : _GEN_42; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_44 = 8'h2c == io_in_0 ? 8'h58 : _GEN_43; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_45 = 8'h2d == io_in_0 ? 8'h5a : _GEN_44; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_46 = 8'h2e == io_in_0 ? 8'h5c : _GEN_45; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_47 = 8'h2f == io_in_0 ? 8'h5e : _GEN_46; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_48 = 8'h30 == io_in_0 ? 8'h60 : _GEN_47; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_49 = 8'h31 == io_in_0 ? 8'h62 : _GEN_48; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_50 = 8'h32 == io_in_0 ? 8'h64 : _GEN_49; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_51 = 8'h33 == io_in_0 ? 8'h66 : _GEN_50; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_52 = 8'h34 == io_in_0 ? 8'h68 : _GEN_51; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_53 = 8'h35 == io_in_0 ? 8'h6a : _GEN_52; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_54 = 8'h36 == io_in_0 ? 8'h6c : _GEN_53; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_55 = 8'h37 == io_in_0 ? 8'h6e : _GEN_54; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_56 = 8'h38 == io_in_0 ? 8'h70 : _GEN_55; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_57 = 8'h39 == io_in_0 ? 8'h72 : _GEN_56; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_58 = 8'h3a == io_in_0 ? 8'h74 : _GEN_57; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_59 = 8'h3b == io_in_0 ? 8'h76 : _GEN_58; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_60 = 8'h3c == io_in_0 ? 8'h78 : _GEN_59; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_61 = 8'h3d == io_in_0 ? 8'h7a : _GEN_60; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_62 = 8'h3e == io_in_0 ? 8'h7c : _GEN_61; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_63 = 8'h3f == io_in_0 ? 8'h7e : _GEN_62; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_64 = 8'h40 == io_in_0 ? 8'h80 : _GEN_63; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_65 = 8'h41 == io_in_0 ? 8'h82 : _GEN_64; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_66 = 8'h42 == io_in_0 ? 8'h84 : _GEN_65; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_67 = 8'h43 == io_in_0 ? 8'h86 : _GEN_66; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_68 = 8'h44 == io_in_0 ? 8'h88 : _GEN_67; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_69 = 8'h45 == io_in_0 ? 8'h8a : _GEN_68; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_70 = 8'h46 == io_in_0 ? 8'h8c : _GEN_69; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_71 = 8'h47 == io_in_0 ? 8'h8e : _GEN_70; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_72 = 8'h48 == io_in_0 ? 8'h90 : _GEN_71; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_73 = 8'h49 == io_in_0 ? 8'h92 : _GEN_72; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_74 = 8'h4a == io_in_0 ? 8'h94 : _GEN_73; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_75 = 8'h4b == io_in_0 ? 8'h96 : _GEN_74; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_76 = 8'h4c == io_in_0 ? 8'h98 : _GEN_75; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_77 = 8'h4d == io_in_0 ? 8'h9a : _GEN_76; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_78 = 8'h4e == io_in_0 ? 8'h9c : _GEN_77; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_79 = 8'h4f == io_in_0 ? 8'h9e : _GEN_78; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_80 = 8'h50 == io_in_0 ? 8'ha0 : _GEN_79; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_81 = 8'h51 == io_in_0 ? 8'ha2 : _GEN_80; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_82 = 8'h52 == io_in_0 ? 8'ha4 : _GEN_81; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_83 = 8'h53 == io_in_0 ? 8'ha6 : _GEN_82; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_84 = 8'h54 == io_in_0 ? 8'ha8 : _GEN_83; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_85 = 8'h55 == io_in_0 ? 8'haa : _GEN_84; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_86 = 8'h56 == io_in_0 ? 8'hac : _GEN_85; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_87 = 8'h57 == io_in_0 ? 8'hae : _GEN_86; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_88 = 8'h58 == io_in_0 ? 8'hb0 : _GEN_87; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_89 = 8'h59 == io_in_0 ? 8'hb2 : _GEN_88; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_90 = 8'h5a == io_in_0 ? 8'hb4 : _GEN_89; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_91 = 8'h5b == io_in_0 ? 8'hb6 : _GEN_90; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_92 = 8'h5c == io_in_0 ? 8'hb8 : _GEN_91; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_93 = 8'h5d == io_in_0 ? 8'hba : _GEN_92; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_94 = 8'h5e == io_in_0 ? 8'hbc : _GEN_93; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_95 = 8'h5f == io_in_0 ? 8'hbe : _GEN_94; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_96 = 8'h60 == io_in_0 ? 8'hc0 : _GEN_95; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_97 = 8'h61 == io_in_0 ? 8'hc2 : _GEN_96; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_98 = 8'h62 == io_in_0 ? 8'hc4 : _GEN_97; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_99 = 8'h63 == io_in_0 ? 8'hc6 : _GEN_98; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_100 = 8'h64 == io_in_0 ? 8'hc8 : _GEN_99; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_101 = 8'h65 == io_in_0 ? 8'hca : _GEN_100; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_102 = 8'h66 == io_in_0 ? 8'hcc : _GEN_101; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_103 = 8'h67 == io_in_0 ? 8'hce : _GEN_102; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_104 = 8'h68 == io_in_0 ? 8'hd0 : _GEN_103; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_105 = 8'h69 == io_in_0 ? 8'hd2 : _GEN_104; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_106 = 8'h6a == io_in_0 ? 8'hd4 : _GEN_105; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_107 = 8'h6b == io_in_0 ? 8'hd6 : _GEN_106; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_108 = 8'h6c == io_in_0 ? 8'hd8 : _GEN_107; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_109 = 8'h6d == io_in_0 ? 8'hda : _GEN_108; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_110 = 8'h6e == io_in_0 ? 8'hdc : _GEN_109; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_111 = 8'h6f == io_in_0 ? 8'hde : _GEN_110; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_112 = 8'h70 == io_in_0 ? 8'he0 : _GEN_111; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_113 = 8'h71 == io_in_0 ? 8'he2 : _GEN_112; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_114 = 8'h72 == io_in_0 ? 8'he4 : _GEN_113; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_115 = 8'h73 == io_in_0 ? 8'he6 : _GEN_114; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_116 = 8'h74 == io_in_0 ? 8'he8 : _GEN_115; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_117 = 8'h75 == io_in_0 ? 8'hea : _GEN_116; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_118 = 8'h76 == io_in_0 ? 8'hec : _GEN_117; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_119 = 8'h77 == io_in_0 ? 8'hee : _GEN_118; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_120 = 8'h78 == io_in_0 ? 8'hf0 : _GEN_119; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_121 = 8'h79 == io_in_0 ? 8'hf2 : _GEN_120; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_122 = 8'h7a == io_in_0 ? 8'hf4 : _GEN_121; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_123 = 8'h7b == io_in_0 ? 8'hf6 : _GEN_122; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_124 = 8'h7c == io_in_0 ? 8'hf8 : _GEN_123; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_125 = 8'h7d == io_in_0 ? 8'hfa : _GEN_124; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_126 = 8'h7e == io_in_0 ? 8'hfc : _GEN_125; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_127 = 8'h7f == io_in_0 ? 8'hfe : _GEN_126; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_128 = 8'h80 == io_in_0 ? 8'h1b : _GEN_127; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_129 = 8'h81 == io_in_0 ? 8'h19 : _GEN_128; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_130 = 8'h82 == io_in_0 ? 8'h1f : _GEN_129; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_131 = 8'h83 == io_in_0 ? 8'h1d : _GEN_130; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_132 = 8'h84 == io_in_0 ? 8'h13 : _GEN_131; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_133 = 8'h85 == io_in_0 ? 8'h11 : _GEN_132; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_134 = 8'h86 == io_in_0 ? 8'h17 : _GEN_133; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_135 = 8'h87 == io_in_0 ? 8'h15 : _GEN_134; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_136 = 8'h88 == io_in_0 ? 8'hb : _GEN_135; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_137 = 8'h89 == io_in_0 ? 8'h9 : _GEN_136; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_138 = 8'h8a == io_in_0 ? 8'hf : _GEN_137; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_139 = 8'h8b == io_in_0 ? 8'hd : _GEN_138; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_140 = 8'h8c == io_in_0 ? 8'h3 : _GEN_139; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_141 = 8'h8d == io_in_0 ? 8'h1 : _GEN_140; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_142 = 8'h8e == io_in_0 ? 8'h7 : _GEN_141; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_143 = 8'h8f == io_in_0 ? 8'h5 : _GEN_142; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_144 = 8'h90 == io_in_0 ? 8'h3b : _GEN_143; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_145 = 8'h91 == io_in_0 ? 8'h39 : _GEN_144; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_146 = 8'h92 == io_in_0 ? 8'h3f : _GEN_145; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_147 = 8'h93 == io_in_0 ? 8'h3d : _GEN_146; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_148 = 8'h94 == io_in_0 ? 8'h33 : _GEN_147; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_149 = 8'h95 == io_in_0 ? 8'h31 : _GEN_148; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_150 = 8'h96 == io_in_0 ? 8'h37 : _GEN_149; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_151 = 8'h97 == io_in_0 ? 8'h35 : _GEN_150; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_152 = 8'h98 == io_in_0 ? 8'h2b : _GEN_151; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_153 = 8'h99 == io_in_0 ? 8'h29 : _GEN_152; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_154 = 8'h9a == io_in_0 ? 8'h2f : _GEN_153; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_155 = 8'h9b == io_in_0 ? 8'h2d : _GEN_154; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_156 = 8'h9c == io_in_0 ? 8'h23 : _GEN_155; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_157 = 8'h9d == io_in_0 ? 8'h21 : _GEN_156; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_158 = 8'h9e == io_in_0 ? 8'h27 : _GEN_157; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_159 = 8'h9f == io_in_0 ? 8'h25 : _GEN_158; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_160 = 8'ha0 == io_in_0 ? 8'h5b : _GEN_159; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_161 = 8'ha1 == io_in_0 ? 8'h59 : _GEN_160; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_162 = 8'ha2 == io_in_0 ? 8'h5f : _GEN_161; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_163 = 8'ha3 == io_in_0 ? 8'h5d : _GEN_162; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_164 = 8'ha4 == io_in_0 ? 8'h53 : _GEN_163; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_165 = 8'ha5 == io_in_0 ? 8'h51 : _GEN_164; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_166 = 8'ha6 == io_in_0 ? 8'h57 : _GEN_165; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_167 = 8'ha7 == io_in_0 ? 8'h55 : _GEN_166; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_168 = 8'ha8 == io_in_0 ? 8'h4b : _GEN_167; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_169 = 8'ha9 == io_in_0 ? 8'h49 : _GEN_168; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_170 = 8'haa == io_in_0 ? 8'h4f : _GEN_169; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_171 = 8'hab == io_in_0 ? 8'h4d : _GEN_170; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_172 = 8'hac == io_in_0 ? 8'h43 : _GEN_171; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_173 = 8'had == io_in_0 ? 8'h41 : _GEN_172; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_174 = 8'hae == io_in_0 ? 8'h47 : _GEN_173; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_175 = 8'haf == io_in_0 ? 8'h45 : _GEN_174; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_176 = 8'hb0 == io_in_0 ? 8'h7b : _GEN_175; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_177 = 8'hb1 == io_in_0 ? 8'h79 : _GEN_176; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_178 = 8'hb2 == io_in_0 ? 8'h7f : _GEN_177; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_179 = 8'hb3 == io_in_0 ? 8'h7d : _GEN_178; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_180 = 8'hb4 == io_in_0 ? 8'h73 : _GEN_179; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_181 = 8'hb5 == io_in_0 ? 8'h71 : _GEN_180; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_182 = 8'hb6 == io_in_0 ? 8'h77 : _GEN_181; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_183 = 8'hb7 == io_in_0 ? 8'h75 : _GEN_182; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_184 = 8'hb8 == io_in_0 ? 8'h6b : _GEN_183; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_185 = 8'hb9 == io_in_0 ? 8'h69 : _GEN_184; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_186 = 8'hba == io_in_0 ? 8'h6f : _GEN_185; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_187 = 8'hbb == io_in_0 ? 8'h6d : _GEN_186; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_188 = 8'hbc == io_in_0 ? 8'h63 : _GEN_187; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_189 = 8'hbd == io_in_0 ? 8'h61 : _GEN_188; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_190 = 8'hbe == io_in_0 ? 8'h67 : _GEN_189; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_191 = 8'hbf == io_in_0 ? 8'h65 : _GEN_190; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_192 = 8'hc0 == io_in_0 ? 8'h9b : _GEN_191; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_193 = 8'hc1 == io_in_0 ? 8'h99 : _GEN_192; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_194 = 8'hc2 == io_in_0 ? 8'h9f : _GEN_193; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_195 = 8'hc3 == io_in_0 ? 8'h9d : _GEN_194; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_196 = 8'hc4 == io_in_0 ? 8'h93 : _GEN_195; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_197 = 8'hc5 == io_in_0 ? 8'h91 : _GEN_196; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_198 = 8'hc6 == io_in_0 ? 8'h97 : _GEN_197; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_199 = 8'hc7 == io_in_0 ? 8'h95 : _GEN_198; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_200 = 8'hc8 == io_in_0 ? 8'h8b : _GEN_199; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_201 = 8'hc9 == io_in_0 ? 8'h89 : _GEN_200; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_202 = 8'hca == io_in_0 ? 8'h8f : _GEN_201; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_203 = 8'hcb == io_in_0 ? 8'h8d : _GEN_202; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_204 = 8'hcc == io_in_0 ? 8'h83 : _GEN_203; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_205 = 8'hcd == io_in_0 ? 8'h81 : _GEN_204; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_206 = 8'hce == io_in_0 ? 8'h87 : _GEN_205; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_207 = 8'hcf == io_in_0 ? 8'h85 : _GEN_206; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_208 = 8'hd0 == io_in_0 ? 8'hbb : _GEN_207; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_209 = 8'hd1 == io_in_0 ? 8'hb9 : _GEN_208; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_210 = 8'hd2 == io_in_0 ? 8'hbf : _GEN_209; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_211 = 8'hd3 == io_in_0 ? 8'hbd : _GEN_210; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_212 = 8'hd4 == io_in_0 ? 8'hb3 : _GEN_211; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_213 = 8'hd5 == io_in_0 ? 8'hb1 : _GEN_212; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_214 = 8'hd6 == io_in_0 ? 8'hb7 : _GEN_213; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_215 = 8'hd7 == io_in_0 ? 8'hb5 : _GEN_214; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_216 = 8'hd8 == io_in_0 ? 8'hab : _GEN_215; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_217 = 8'hd9 == io_in_0 ? 8'ha9 : _GEN_216; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_218 = 8'hda == io_in_0 ? 8'haf : _GEN_217; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_219 = 8'hdb == io_in_0 ? 8'had : _GEN_218; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_220 = 8'hdc == io_in_0 ? 8'ha3 : _GEN_219; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_221 = 8'hdd == io_in_0 ? 8'ha1 : _GEN_220; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_222 = 8'hde == io_in_0 ? 8'ha7 : _GEN_221; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_223 = 8'hdf == io_in_0 ? 8'ha5 : _GEN_222; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_224 = 8'he0 == io_in_0 ? 8'hdb : _GEN_223; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_225 = 8'he1 == io_in_0 ? 8'hd9 : _GEN_224; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_226 = 8'he2 == io_in_0 ? 8'hdf : _GEN_225; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_227 = 8'he3 == io_in_0 ? 8'hdd : _GEN_226; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_228 = 8'he4 == io_in_0 ? 8'hd3 : _GEN_227; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_229 = 8'he5 == io_in_0 ? 8'hd1 : _GEN_228; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_230 = 8'he6 == io_in_0 ? 8'hd7 : _GEN_229; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_231 = 8'he7 == io_in_0 ? 8'hd5 : _GEN_230; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_232 = 8'he8 == io_in_0 ? 8'hcb : _GEN_231; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_233 = 8'he9 == io_in_0 ? 8'hc9 : _GEN_232; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_234 = 8'hea == io_in_0 ? 8'hcf : _GEN_233; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_235 = 8'heb == io_in_0 ? 8'hcd : _GEN_234; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_236 = 8'hec == io_in_0 ? 8'hc3 : _GEN_235; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_237 = 8'hed == io_in_0 ? 8'hc1 : _GEN_236; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_238 = 8'hee == io_in_0 ? 8'hc7 : _GEN_237; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_239 = 8'hef == io_in_0 ? 8'hc5 : _GEN_238; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_240 = 8'hf0 == io_in_0 ? 8'hfb : _GEN_239; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_241 = 8'hf1 == io_in_0 ? 8'hf9 : _GEN_240; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_242 = 8'hf2 == io_in_0 ? 8'hff : _GEN_241; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_243 = 8'hf3 == io_in_0 ? 8'hfd : _GEN_242; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_244 = 8'hf4 == io_in_0 ? 8'hf3 : _GEN_243; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_245 = 8'hf5 == io_in_0 ? 8'hf1 : _GEN_244; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_246 = 8'hf6 == io_in_0 ? 8'hf7 : _GEN_245; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_247 = 8'hf7 == io_in_0 ? 8'hf5 : _GEN_246; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_248 = 8'hf8 == io_in_0 ? 8'heb : _GEN_247; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_249 = 8'hf9 == io_in_0 ? 8'he9 : _GEN_248; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_250 = 8'hfa == io_in_0 ? 8'hef : _GEN_249; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_251 = 8'hfb == io_in_0 ? 8'hed : _GEN_250; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_252 = 8'hfc == io_in_0 ? 8'he3 : _GEN_251; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_253 = 8'hfd == io_in_0 ? 8'he1 : _GEN_252; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_254 = 8'hfe == io_in_0 ? 8'he7 : _GEN_253; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_255 = 8'hff == io_in_0 ? 8'he5 : _GEN_254; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_257 = 8'h1 == io_in_1 ? 8'h2 : 8'h0; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_258 = 8'h2 == io_in_1 ? 8'h4 : _GEN_257; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_259 = 8'h3 == io_in_1 ? 8'h6 : _GEN_258; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_260 = 8'h4 == io_in_1 ? 8'h8 : _GEN_259; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_261 = 8'h5 == io_in_1 ? 8'ha : _GEN_260; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_262 = 8'h6 == io_in_1 ? 8'hc : _GEN_261; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_263 = 8'h7 == io_in_1 ? 8'he : _GEN_262; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_264 = 8'h8 == io_in_1 ? 8'h10 : _GEN_263; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_265 = 8'h9 == io_in_1 ? 8'h12 : _GEN_264; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_266 = 8'ha == io_in_1 ? 8'h14 : _GEN_265; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_267 = 8'hb == io_in_1 ? 8'h16 : _GEN_266; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_268 = 8'hc == io_in_1 ? 8'h18 : _GEN_267; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_269 = 8'hd == io_in_1 ? 8'h1a : _GEN_268; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_270 = 8'he == io_in_1 ? 8'h1c : _GEN_269; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_271 = 8'hf == io_in_1 ? 8'h1e : _GEN_270; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_272 = 8'h10 == io_in_1 ? 8'h20 : _GEN_271; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_273 = 8'h11 == io_in_1 ? 8'h22 : _GEN_272; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_274 = 8'h12 == io_in_1 ? 8'h24 : _GEN_273; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_275 = 8'h13 == io_in_1 ? 8'h26 : _GEN_274; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_276 = 8'h14 == io_in_1 ? 8'h28 : _GEN_275; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_277 = 8'h15 == io_in_1 ? 8'h2a : _GEN_276; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_278 = 8'h16 == io_in_1 ? 8'h2c : _GEN_277; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_279 = 8'h17 == io_in_1 ? 8'h2e : _GEN_278; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_280 = 8'h18 == io_in_1 ? 8'h30 : _GEN_279; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_281 = 8'h19 == io_in_1 ? 8'h32 : _GEN_280; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_282 = 8'h1a == io_in_1 ? 8'h34 : _GEN_281; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_283 = 8'h1b == io_in_1 ? 8'h36 : _GEN_282; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_284 = 8'h1c == io_in_1 ? 8'h38 : _GEN_283; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_285 = 8'h1d == io_in_1 ? 8'h3a : _GEN_284; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_286 = 8'h1e == io_in_1 ? 8'h3c : _GEN_285; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_287 = 8'h1f == io_in_1 ? 8'h3e : _GEN_286; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_288 = 8'h20 == io_in_1 ? 8'h40 : _GEN_287; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_289 = 8'h21 == io_in_1 ? 8'h42 : _GEN_288; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_290 = 8'h22 == io_in_1 ? 8'h44 : _GEN_289; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_291 = 8'h23 == io_in_1 ? 8'h46 : _GEN_290; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_292 = 8'h24 == io_in_1 ? 8'h48 : _GEN_291; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_293 = 8'h25 == io_in_1 ? 8'h4a : _GEN_292; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_294 = 8'h26 == io_in_1 ? 8'h4c : _GEN_293; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_295 = 8'h27 == io_in_1 ? 8'h4e : _GEN_294; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_296 = 8'h28 == io_in_1 ? 8'h50 : _GEN_295; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_297 = 8'h29 == io_in_1 ? 8'h52 : _GEN_296; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_298 = 8'h2a == io_in_1 ? 8'h54 : _GEN_297; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_299 = 8'h2b == io_in_1 ? 8'h56 : _GEN_298; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_300 = 8'h2c == io_in_1 ? 8'h58 : _GEN_299; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_301 = 8'h2d == io_in_1 ? 8'h5a : _GEN_300; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_302 = 8'h2e == io_in_1 ? 8'h5c : _GEN_301; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_303 = 8'h2f == io_in_1 ? 8'h5e : _GEN_302; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_304 = 8'h30 == io_in_1 ? 8'h60 : _GEN_303; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_305 = 8'h31 == io_in_1 ? 8'h62 : _GEN_304; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_306 = 8'h32 == io_in_1 ? 8'h64 : _GEN_305; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_307 = 8'h33 == io_in_1 ? 8'h66 : _GEN_306; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_308 = 8'h34 == io_in_1 ? 8'h68 : _GEN_307; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_309 = 8'h35 == io_in_1 ? 8'h6a : _GEN_308; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_310 = 8'h36 == io_in_1 ? 8'h6c : _GEN_309; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_311 = 8'h37 == io_in_1 ? 8'h6e : _GEN_310; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_312 = 8'h38 == io_in_1 ? 8'h70 : _GEN_311; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_313 = 8'h39 == io_in_1 ? 8'h72 : _GEN_312; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_314 = 8'h3a == io_in_1 ? 8'h74 : _GEN_313; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_315 = 8'h3b == io_in_1 ? 8'h76 : _GEN_314; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_316 = 8'h3c == io_in_1 ? 8'h78 : _GEN_315; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_317 = 8'h3d == io_in_1 ? 8'h7a : _GEN_316; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_318 = 8'h3e == io_in_1 ? 8'h7c : _GEN_317; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_319 = 8'h3f == io_in_1 ? 8'h7e : _GEN_318; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_320 = 8'h40 == io_in_1 ? 8'h80 : _GEN_319; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_321 = 8'h41 == io_in_1 ? 8'h82 : _GEN_320; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_322 = 8'h42 == io_in_1 ? 8'h84 : _GEN_321; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_323 = 8'h43 == io_in_1 ? 8'h86 : _GEN_322; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_324 = 8'h44 == io_in_1 ? 8'h88 : _GEN_323; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_325 = 8'h45 == io_in_1 ? 8'h8a : _GEN_324; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_326 = 8'h46 == io_in_1 ? 8'h8c : _GEN_325; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_327 = 8'h47 == io_in_1 ? 8'h8e : _GEN_326; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_328 = 8'h48 == io_in_1 ? 8'h90 : _GEN_327; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_329 = 8'h49 == io_in_1 ? 8'h92 : _GEN_328; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_330 = 8'h4a == io_in_1 ? 8'h94 : _GEN_329; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_331 = 8'h4b == io_in_1 ? 8'h96 : _GEN_330; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_332 = 8'h4c == io_in_1 ? 8'h98 : _GEN_331; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_333 = 8'h4d == io_in_1 ? 8'h9a : _GEN_332; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_334 = 8'h4e == io_in_1 ? 8'h9c : _GEN_333; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_335 = 8'h4f == io_in_1 ? 8'h9e : _GEN_334; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_336 = 8'h50 == io_in_1 ? 8'ha0 : _GEN_335; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_337 = 8'h51 == io_in_1 ? 8'ha2 : _GEN_336; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_338 = 8'h52 == io_in_1 ? 8'ha4 : _GEN_337; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_339 = 8'h53 == io_in_1 ? 8'ha6 : _GEN_338; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_340 = 8'h54 == io_in_1 ? 8'ha8 : _GEN_339; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_341 = 8'h55 == io_in_1 ? 8'haa : _GEN_340; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_342 = 8'h56 == io_in_1 ? 8'hac : _GEN_341; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_343 = 8'h57 == io_in_1 ? 8'hae : _GEN_342; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_344 = 8'h58 == io_in_1 ? 8'hb0 : _GEN_343; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_345 = 8'h59 == io_in_1 ? 8'hb2 : _GEN_344; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_346 = 8'h5a == io_in_1 ? 8'hb4 : _GEN_345; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_347 = 8'h5b == io_in_1 ? 8'hb6 : _GEN_346; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_348 = 8'h5c == io_in_1 ? 8'hb8 : _GEN_347; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_349 = 8'h5d == io_in_1 ? 8'hba : _GEN_348; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_350 = 8'h5e == io_in_1 ? 8'hbc : _GEN_349; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_351 = 8'h5f == io_in_1 ? 8'hbe : _GEN_350; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_352 = 8'h60 == io_in_1 ? 8'hc0 : _GEN_351; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_353 = 8'h61 == io_in_1 ? 8'hc2 : _GEN_352; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_354 = 8'h62 == io_in_1 ? 8'hc4 : _GEN_353; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_355 = 8'h63 == io_in_1 ? 8'hc6 : _GEN_354; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_356 = 8'h64 == io_in_1 ? 8'hc8 : _GEN_355; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_357 = 8'h65 == io_in_1 ? 8'hca : _GEN_356; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_358 = 8'h66 == io_in_1 ? 8'hcc : _GEN_357; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_359 = 8'h67 == io_in_1 ? 8'hce : _GEN_358; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_360 = 8'h68 == io_in_1 ? 8'hd0 : _GEN_359; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_361 = 8'h69 == io_in_1 ? 8'hd2 : _GEN_360; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_362 = 8'h6a == io_in_1 ? 8'hd4 : _GEN_361; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_363 = 8'h6b == io_in_1 ? 8'hd6 : _GEN_362; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_364 = 8'h6c == io_in_1 ? 8'hd8 : _GEN_363; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_365 = 8'h6d == io_in_1 ? 8'hda : _GEN_364; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_366 = 8'h6e == io_in_1 ? 8'hdc : _GEN_365; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_367 = 8'h6f == io_in_1 ? 8'hde : _GEN_366; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_368 = 8'h70 == io_in_1 ? 8'he0 : _GEN_367; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_369 = 8'h71 == io_in_1 ? 8'he2 : _GEN_368; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_370 = 8'h72 == io_in_1 ? 8'he4 : _GEN_369; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_371 = 8'h73 == io_in_1 ? 8'he6 : _GEN_370; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_372 = 8'h74 == io_in_1 ? 8'he8 : _GEN_371; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_373 = 8'h75 == io_in_1 ? 8'hea : _GEN_372; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_374 = 8'h76 == io_in_1 ? 8'hec : _GEN_373; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_375 = 8'h77 == io_in_1 ? 8'hee : _GEN_374; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_376 = 8'h78 == io_in_1 ? 8'hf0 : _GEN_375; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_377 = 8'h79 == io_in_1 ? 8'hf2 : _GEN_376; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_378 = 8'h7a == io_in_1 ? 8'hf4 : _GEN_377; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_379 = 8'h7b == io_in_1 ? 8'hf6 : _GEN_378; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_380 = 8'h7c == io_in_1 ? 8'hf8 : _GEN_379; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_381 = 8'h7d == io_in_1 ? 8'hfa : _GEN_380; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_382 = 8'h7e == io_in_1 ? 8'hfc : _GEN_381; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_383 = 8'h7f == io_in_1 ? 8'hfe : _GEN_382; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_384 = 8'h80 == io_in_1 ? 8'h1b : _GEN_383; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_385 = 8'h81 == io_in_1 ? 8'h19 : _GEN_384; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_386 = 8'h82 == io_in_1 ? 8'h1f : _GEN_385; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_387 = 8'h83 == io_in_1 ? 8'h1d : _GEN_386; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_388 = 8'h84 == io_in_1 ? 8'h13 : _GEN_387; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_389 = 8'h85 == io_in_1 ? 8'h11 : _GEN_388; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_390 = 8'h86 == io_in_1 ? 8'h17 : _GEN_389; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_391 = 8'h87 == io_in_1 ? 8'h15 : _GEN_390; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_392 = 8'h88 == io_in_1 ? 8'hb : _GEN_391; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_393 = 8'h89 == io_in_1 ? 8'h9 : _GEN_392; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_394 = 8'h8a == io_in_1 ? 8'hf : _GEN_393; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_395 = 8'h8b == io_in_1 ? 8'hd : _GEN_394; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_396 = 8'h8c == io_in_1 ? 8'h3 : _GEN_395; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_397 = 8'h8d == io_in_1 ? 8'h1 : _GEN_396; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_398 = 8'h8e == io_in_1 ? 8'h7 : _GEN_397; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_399 = 8'h8f == io_in_1 ? 8'h5 : _GEN_398; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_400 = 8'h90 == io_in_1 ? 8'h3b : _GEN_399; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_401 = 8'h91 == io_in_1 ? 8'h39 : _GEN_400; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_402 = 8'h92 == io_in_1 ? 8'h3f : _GEN_401; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_403 = 8'h93 == io_in_1 ? 8'h3d : _GEN_402; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_404 = 8'h94 == io_in_1 ? 8'h33 : _GEN_403; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_405 = 8'h95 == io_in_1 ? 8'h31 : _GEN_404; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_406 = 8'h96 == io_in_1 ? 8'h37 : _GEN_405; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_407 = 8'h97 == io_in_1 ? 8'h35 : _GEN_406; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_408 = 8'h98 == io_in_1 ? 8'h2b : _GEN_407; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_409 = 8'h99 == io_in_1 ? 8'h29 : _GEN_408; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_410 = 8'h9a == io_in_1 ? 8'h2f : _GEN_409; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_411 = 8'h9b == io_in_1 ? 8'h2d : _GEN_410; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_412 = 8'h9c == io_in_1 ? 8'h23 : _GEN_411; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_413 = 8'h9d == io_in_1 ? 8'h21 : _GEN_412; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_414 = 8'h9e == io_in_1 ? 8'h27 : _GEN_413; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_415 = 8'h9f == io_in_1 ? 8'h25 : _GEN_414; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_416 = 8'ha0 == io_in_1 ? 8'h5b : _GEN_415; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_417 = 8'ha1 == io_in_1 ? 8'h59 : _GEN_416; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_418 = 8'ha2 == io_in_1 ? 8'h5f : _GEN_417; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_419 = 8'ha3 == io_in_1 ? 8'h5d : _GEN_418; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_420 = 8'ha4 == io_in_1 ? 8'h53 : _GEN_419; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_421 = 8'ha5 == io_in_1 ? 8'h51 : _GEN_420; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_422 = 8'ha6 == io_in_1 ? 8'h57 : _GEN_421; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_423 = 8'ha7 == io_in_1 ? 8'h55 : _GEN_422; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_424 = 8'ha8 == io_in_1 ? 8'h4b : _GEN_423; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_425 = 8'ha9 == io_in_1 ? 8'h49 : _GEN_424; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_426 = 8'haa == io_in_1 ? 8'h4f : _GEN_425; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_427 = 8'hab == io_in_1 ? 8'h4d : _GEN_426; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_428 = 8'hac == io_in_1 ? 8'h43 : _GEN_427; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_429 = 8'had == io_in_1 ? 8'h41 : _GEN_428; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_430 = 8'hae == io_in_1 ? 8'h47 : _GEN_429; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_431 = 8'haf == io_in_1 ? 8'h45 : _GEN_430; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_432 = 8'hb0 == io_in_1 ? 8'h7b : _GEN_431; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_433 = 8'hb1 == io_in_1 ? 8'h79 : _GEN_432; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_434 = 8'hb2 == io_in_1 ? 8'h7f : _GEN_433; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_435 = 8'hb3 == io_in_1 ? 8'h7d : _GEN_434; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_436 = 8'hb4 == io_in_1 ? 8'h73 : _GEN_435; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_437 = 8'hb5 == io_in_1 ? 8'h71 : _GEN_436; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_438 = 8'hb6 == io_in_1 ? 8'h77 : _GEN_437; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_439 = 8'hb7 == io_in_1 ? 8'h75 : _GEN_438; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_440 = 8'hb8 == io_in_1 ? 8'h6b : _GEN_439; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_441 = 8'hb9 == io_in_1 ? 8'h69 : _GEN_440; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_442 = 8'hba == io_in_1 ? 8'h6f : _GEN_441; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_443 = 8'hbb == io_in_1 ? 8'h6d : _GEN_442; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_444 = 8'hbc == io_in_1 ? 8'h63 : _GEN_443; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_445 = 8'hbd == io_in_1 ? 8'h61 : _GEN_444; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_446 = 8'hbe == io_in_1 ? 8'h67 : _GEN_445; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_447 = 8'hbf == io_in_1 ? 8'h65 : _GEN_446; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_448 = 8'hc0 == io_in_1 ? 8'h9b : _GEN_447; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_449 = 8'hc1 == io_in_1 ? 8'h99 : _GEN_448; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_450 = 8'hc2 == io_in_1 ? 8'h9f : _GEN_449; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_451 = 8'hc3 == io_in_1 ? 8'h9d : _GEN_450; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_452 = 8'hc4 == io_in_1 ? 8'h93 : _GEN_451; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_453 = 8'hc5 == io_in_1 ? 8'h91 : _GEN_452; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_454 = 8'hc6 == io_in_1 ? 8'h97 : _GEN_453; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_455 = 8'hc7 == io_in_1 ? 8'h95 : _GEN_454; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_456 = 8'hc8 == io_in_1 ? 8'h8b : _GEN_455; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_457 = 8'hc9 == io_in_1 ? 8'h89 : _GEN_456; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_458 = 8'hca == io_in_1 ? 8'h8f : _GEN_457; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_459 = 8'hcb == io_in_1 ? 8'h8d : _GEN_458; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_460 = 8'hcc == io_in_1 ? 8'h83 : _GEN_459; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_461 = 8'hcd == io_in_1 ? 8'h81 : _GEN_460; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_462 = 8'hce == io_in_1 ? 8'h87 : _GEN_461; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_463 = 8'hcf == io_in_1 ? 8'h85 : _GEN_462; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_464 = 8'hd0 == io_in_1 ? 8'hbb : _GEN_463; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_465 = 8'hd1 == io_in_1 ? 8'hb9 : _GEN_464; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_466 = 8'hd2 == io_in_1 ? 8'hbf : _GEN_465; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_467 = 8'hd3 == io_in_1 ? 8'hbd : _GEN_466; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_468 = 8'hd4 == io_in_1 ? 8'hb3 : _GEN_467; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_469 = 8'hd5 == io_in_1 ? 8'hb1 : _GEN_468; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_470 = 8'hd6 == io_in_1 ? 8'hb7 : _GEN_469; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_471 = 8'hd7 == io_in_1 ? 8'hb5 : _GEN_470; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_472 = 8'hd8 == io_in_1 ? 8'hab : _GEN_471; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_473 = 8'hd9 == io_in_1 ? 8'ha9 : _GEN_472; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_474 = 8'hda == io_in_1 ? 8'haf : _GEN_473; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_475 = 8'hdb == io_in_1 ? 8'had : _GEN_474; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_476 = 8'hdc == io_in_1 ? 8'ha3 : _GEN_475; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_477 = 8'hdd == io_in_1 ? 8'ha1 : _GEN_476; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_478 = 8'hde == io_in_1 ? 8'ha7 : _GEN_477; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_479 = 8'hdf == io_in_1 ? 8'ha5 : _GEN_478; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_480 = 8'he0 == io_in_1 ? 8'hdb : _GEN_479; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_481 = 8'he1 == io_in_1 ? 8'hd9 : _GEN_480; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_482 = 8'he2 == io_in_1 ? 8'hdf : _GEN_481; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_483 = 8'he3 == io_in_1 ? 8'hdd : _GEN_482; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_484 = 8'he4 == io_in_1 ? 8'hd3 : _GEN_483; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_485 = 8'he5 == io_in_1 ? 8'hd1 : _GEN_484; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_486 = 8'he6 == io_in_1 ? 8'hd7 : _GEN_485; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_487 = 8'he7 == io_in_1 ? 8'hd5 : _GEN_486; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_488 = 8'he8 == io_in_1 ? 8'hcb : _GEN_487; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_489 = 8'he9 == io_in_1 ? 8'hc9 : _GEN_488; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_490 = 8'hea == io_in_1 ? 8'hcf : _GEN_489; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_491 = 8'heb == io_in_1 ? 8'hcd : _GEN_490; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_492 = 8'hec == io_in_1 ? 8'hc3 : _GEN_491; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_493 = 8'hed == io_in_1 ? 8'hc1 : _GEN_492; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_494 = 8'hee == io_in_1 ? 8'hc7 : _GEN_493; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_495 = 8'hef == io_in_1 ? 8'hc5 : _GEN_494; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_496 = 8'hf0 == io_in_1 ? 8'hfb : _GEN_495; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_497 = 8'hf1 == io_in_1 ? 8'hf9 : _GEN_496; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_498 = 8'hf2 == io_in_1 ? 8'hff : _GEN_497; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_499 = 8'hf3 == io_in_1 ? 8'hfd : _GEN_498; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_500 = 8'hf4 == io_in_1 ? 8'hf3 : _GEN_499; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_501 = 8'hf5 == io_in_1 ? 8'hf1 : _GEN_500; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_502 = 8'hf6 == io_in_1 ? 8'hf7 : _GEN_501; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_503 = 8'hf7 == io_in_1 ? 8'hf5 : _GEN_502; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_504 = 8'hf8 == io_in_1 ? 8'heb : _GEN_503; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_505 = 8'hf9 == io_in_1 ? 8'he9 : _GEN_504; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_506 = 8'hfa == io_in_1 ? 8'hef : _GEN_505; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_507 = 8'hfb == io_in_1 ? 8'hed : _GEN_506; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_508 = 8'hfc == io_in_1 ? 8'he3 : _GEN_507; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_509 = 8'hfd == io_in_1 ? 8'he1 : _GEN_508; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_510 = 8'hfe == io_in_1 ? 8'he7 : _GEN_509; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _GEN_511 = 8'hff == io_in_1 ? 8'he5 : _GEN_510; // @[AES_EncryptionFSM.scala 296:31 AES_EncryptionFSM.scala 296:31]
  wire [7:0] _T = _GEN_255 ^ _GEN_511; // @[AES_EncryptionFSM.scala 296:31]
  wire [7:0] _T_1 = _T ^ io_in_1; // @[AES_EncryptionFSM.scala 296:48]
  wire [7:0] _T_2 = _T_1 ^ io_in_2; // @[AES_EncryptionFSM.scala 296:59]
  wire [7:0] _T_4 = io_in_0 ^ _GEN_511; // @[AES_EncryptionFSM.scala 297:25]
  wire [7:0] _GEN_513 = 8'h1 == io_in_2 ? 8'h2 : 8'h0; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_514 = 8'h2 == io_in_2 ? 8'h4 : _GEN_513; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_515 = 8'h3 == io_in_2 ? 8'h6 : _GEN_514; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_516 = 8'h4 == io_in_2 ? 8'h8 : _GEN_515; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_517 = 8'h5 == io_in_2 ? 8'ha : _GEN_516; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_518 = 8'h6 == io_in_2 ? 8'hc : _GEN_517; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_519 = 8'h7 == io_in_2 ? 8'he : _GEN_518; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_520 = 8'h8 == io_in_2 ? 8'h10 : _GEN_519; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_521 = 8'h9 == io_in_2 ? 8'h12 : _GEN_520; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_522 = 8'ha == io_in_2 ? 8'h14 : _GEN_521; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_523 = 8'hb == io_in_2 ? 8'h16 : _GEN_522; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_524 = 8'hc == io_in_2 ? 8'h18 : _GEN_523; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_525 = 8'hd == io_in_2 ? 8'h1a : _GEN_524; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_526 = 8'he == io_in_2 ? 8'h1c : _GEN_525; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_527 = 8'hf == io_in_2 ? 8'h1e : _GEN_526; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_528 = 8'h10 == io_in_2 ? 8'h20 : _GEN_527; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_529 = 8'h11 == io_in_2 ? 8'h22 : _GEN_528; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_530 = 8'h12 == io_in_2 ? 8'h24 : _GEN_529; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_531 = 8'h13 == io_in_2 ? 8'h26 : _GEN_530; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_532 = 8'h14 == io_in_2 ? 8'h28 : _GEN_531; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_533 = 8'h15 == io_in_2 ? 8'h2a : _GEN_532; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_534 = 8'h16 == io_in_2 ? 8'h2c : _GEN_533; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_535 = 8'h17 == io_in_2 ? 8'h2e : _GEN_534; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_536 = 8'h18 == io_in_2 ? 8'h30 : _GEN_535; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_537 = 8'h19 == io_in_2 ? 8'h32 : _GEN_536; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_538 = 8'h1a == io_in_2 ? 8'h34 : _GEN_537; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_539 = 8'h1b == io_in_2 ? 8'h36 : _GEN_538; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_540 = 8'h1c == io_in_2 ? 8'h38 : _GEN_539; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_541 = 8'h1d == io_in_2 ? 8'h3a : _GEN_540; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_542 = 8'h1e == io_in_2 ? 8'h3c : _GEN_541; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_543 = 8'h1f == io_in_2 ? 8'h3e : _GEN_542; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_544 = 8'h20 == io_in_2 ? 8'h40 : _GEN_543; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_545 = 8'h21 == io_in_2 ? 8'h42 : _GEN_544; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_546 = 8'h22 == io_in_2 ? 8'h44 : _GEN_545; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_547 = 8'h23 == io_in_2 ? 8'h46 : _GEN_546; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_548 = 8'h24 == io_in_2 ? 8'h48 : _GEN_547; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_549 = 8'h25 == io_in_2 ? 8'h4a : _GEN_548; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_550 = 8'h26 == io_in_2 ? 8'h4c : _GEN_549; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_551 = 8'h27 == io_in_2 ? 8'h4e : _GEN_550; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_552 = 8'h28 == io_in_2 ? 8'h50 : _GEN_551; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_553 = 8'h29 == io_in_2 ? 8'h52 : _GEN_552; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_554 = 8'h2a == io_in_2 ? 8'h54 : _GEN_553; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_555 = 8'h2b == io_in_2 ? 8'h56 : _GEN_554; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_556 = 8'h2c == io_in_2 ? 8'h58 : _GEN_555; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_557 = 8'h2d == io_in_2 ? 8'h5a : _GEN_556; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_558 = 8'h2e == io_in_2 ? 8'h5c : _GEN_557; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_559 = 8'h2f == io_in_2 ? 8'h5e : _GEN_558; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_560 = 8'h30 == io_in_2 ? 8'h60 : _GEN_559; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_561 = 8'h31 == io_in_2 ? 8'h62 : _GEN_560; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_562 = 8'h32 == io_in_2 ? 8'h64 : _GEN_561; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_563 = 8'h33 == io_in_2 ? 8'h66 : _GEN_562; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_564 = 8'h34 == io_in_2 ? 8'h68 : _GEN_563; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_565 = 8'h35 == io_in_2 ? 8'h6a : _GEN_564; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_566 = 8'h36 == io_in_2 ? 8'h6c : _GEN_565; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_567 = 8'h37 == io_in_2 ? 8'h6e : _GEN_566; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_568 = 8'h38 == io_in_2 ? 8'h70 : _GEN_567; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_569 = 8'h39 == io_in_2 ? 8'h72 : _GEN_568; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_570 = 8'h3a == io_in_2 ? 8'h74 : _GEN_569; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_571 = 8'h3b == io_in_2 ? 8'h76 : _GEN_570; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_572 = 8'h3c == io_in_2 ? 8'h78 : _GEN_571; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_573 = 8'h3d == io_in_2 ? 8'h7a : _GEN_572; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_574 = 8'h3e == io_in_2 ? 8'h7c : _GEN_573; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_575 = 8'h3f == io_in_2 ? 8'h7e : _GEN_574; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_576 = 8'h40 == io_in_2 ? 8'h80 : _GEN_575; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_577 = 8'h41 == io_in_2 ? 8'h82 : _GEN_576; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_578 = 8'h42 == io_in_2 ? 8'h84 : _GEN_577; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_579 = 8'h43 == io_in_2 ? 8'h86 : _GEN_578; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_580 = 8'h44 == io_in_2 ? 8'h88 : _GEN_579; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_581 = 8'h45 == io_in_2 ? 8'h8a : _GEN_580; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_582 = 8'h46 == io_in_2 ? 8'h8c : _GEN_581; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_583 = 8'h47 == io_in_2 ? 8'h8e : _GEN_582; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_584 = 8'h48 == io_in_2 ? 8'h90 : _GEN_583; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_585 = 8'h49 == io_in_2 ? 8'h92 : _GEN_584; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_586 = 8'h4a == io_in_2 ? 8'h94 : _GEN_585; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_587 = 8'h4b == io_in_2 ? 8'h96 : _GEN_586; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_588 = 8'h4c == io_in_2 ? 8'h98 : _GEN_587; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_589 = 8'h4d == io_in_2 ? 8'h9a : _GEN_588; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_590 = 8'h4e == io_in_2 ? 8'h9c : _GEN_589; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_591 = 8'h4f == io_in_2 ? 8'h9e : _GEN_590; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_592 = 8'h50 == io_in_2 ? 8'ha0 : _GEN_591; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_593 = 8'h51 == io_in_2 ? 8'ha2 : _GEN_592; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_594 = 8'h52 == io_in_2 ? 8'ha4 : _GEN_593; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_595 = 8'h53 == io_in_2 ? 8'ha6 : _GEN_594; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_596 = 8'h54 == io_in_2 ? 8'ha8 : _GEN_595; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_597 = 8'h55 == io_in_2 ? 8'haa : _GEN_596; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_598 = 8'h56 == io_in_2 ? 8'hac : _GEN_597; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_599 = 8'h57 == io_in_2 ? 8'hae : _GEN_598; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_600 = 8'h58 == io_in_2 ? 8'hb0 : _GEN_599; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_601 = 8'h59 == io_in_2 ? 8'hb2 : _GEN_600; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_602 = 8'h5a == io_in_2 ? 8'hb4 : _GEN_601; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_603 = 8'h5b == io_in_2 ? 8'hb6 : _GEN_602; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_604 = 8'h5c == io_in_2 ? 8'hb8 : _GEN_603; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_605 = 8'h5d == io_in_2 ? 8'hba : _GEN_604; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_606 = 8'h5e == io_in_2 ? 8'hbc : _GEN_605; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_607 = 8'h5f == io_in_2 ? 8'hbe : _GEN_606; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_608 = 8'h60 == io_in_2 ? 8'hc0 : _GEN_607; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_609 = 8'h61 == io_in_2 ? 8'hc2 : _GEN_608; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_610 = 8'h62 == io_in_2 ? 8'hc4 : _GEN_609; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_611 = 8'h63 == io_in_2 ? 8'hc6 : _GEN_610; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_612 = 8'h64 == io_in_2 ? 8'hc8 : _GEN_611; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_613 = 8'h65 == io_in_2 ? 8'hca : _GEN_612; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_614 = 8'h66 == io_in_2 ? 8'hcc : _GEN_613; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_615 = 8'h67 == io_in_2 ? 8'hce : _GEN_614; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_616 = 8'h68 == io_in_2 ? 8'hd0 : _GEN_615; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_617 = 8'h69 == io_in_2 ? 8'hd2 : _GEN_616; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_618 = 8'h6a == io_in_2 ? 8'hd4 : _GEN_617; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_619 = 8'h6b == io_in_2 ? 8'hd6 : _GEN_618; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_620 = 8'h6c == io_in_2 ? 8'hd8 : _GEN_619; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_621 = 8'h6d == io_in_2 ? 8'hda : _GEN_620; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_622 = 8'h6e == io_in_2 ? 8'hdc : _GEN_621; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_623 = 8'h6f == io_in_2 ? 8'hde : _GEN_622; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_624 = 8'h70 == io_in_2 ? 8'he0 : _GEN_623; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_625 = 8'h71 == io_in_2 ? 8'he2 : _GEN_624; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_626 = 8'h72 == io_in_2 ? 8'he4 : _GEN_625; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_627 = 8'h73 == io_in_2 ? 8'he6 : _GEN_626; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_628 = 8'h74 == io_in_2 ? 8'he8 : _GEN_627; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_629 = 8'h75 == io_in_2 ? 8'hea : _GEN_628; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_630 = 8'h76 == io_in_2 ? 8'hec : _GEN_629; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_631 = 8'h77 == io_in_2 ? 8'hee : _GEN_630; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_632 = 8'h78 == io_in_2 ? 8'hf0 : _GEN_631; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_633 = 8'h79 == io_in_2 ? 8'hf2 : _GEN_632; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_634 = 8'h7a == io_in_2 ? 8'hf4 : _GEN_633; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_635 = 8'h7b == io_in_2 ? 8'hf6 : _GEN_634; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_636 = 8'h7c == io_in_2 ? 8'hf8 : _GEN_635; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_637 = 8'h7d == io_in_2 ? 8'hfa : _GEN_636; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_638 = 8'h7e == io_in_2 ? 8'hfc : _GEN_637; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_639 = 8'h7f == io_in_2 ? 8'hfe : _GEN_638; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_640 = 8'h80 == io_in_2 ? 8'h1b : _GEN_639; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_641 = 8'h81 == io_in_2 ? 8'h19 : _GEN_640; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_642 = 8'h82 == io_in_2 ? 8'h1f : _GEN_641; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_643 = 8'h83 == io_in_2 ? 8'h1d : _GEN_642; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_644 = 8'h84 == io_in_2 ? 8'h13 : _GEN_643; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_645 = 8'h85 == io_in_2 ? 8'h11 : _GEN_644; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_646 = 8'h86 == io_in_2 ? 8'h17 : _GEN_645; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_647 = 8'h87 == io_in_2 ? 8'h15 : _GEN_646; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_648 = 8'h88 == io_in_2 ? 8'hb : _GEN_647; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_649 = 8'h89 == io_in_2 ? 8'h9 : _GEN_648; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_650 = 8'h8a == io_in_2 ? 8'hf : _GEN_649; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_651 = 8'h8b == io_in_2 ? 8'hd : _GEN_650; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_652 = 8'h8c == io_in_2 ? 8'h3 : _GEN_651; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_653 = 8'h8d == io_in_2 ? 8'h1 : _GEN_652; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_654 = 8'h8e == io_in_2 ? 8'h7 : _GEN_653; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_655 = 8'h8f == io_in_2 ? 8'h5 : _GEN_654; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_656 = 8'h90 == io_in_2 ? 8'h3b : _GEN_655; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_657 = 8'h91 == io_in_2 ? 8'h39 : _GEN_656; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_658 = 8'h92 == io_in_2 ? 8'h3f : _GEN_657; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_659 = 8'h93 == io_in_2 ? 8'h3d : _GEN_658; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_660 = 8'h94 == io_in_2 ? 8'h33 : _GEN_659; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_661 = 8'h95 == io_in_2 ? 8'h31 : _GEN_660; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_662 = 8'h96 == io_in_2 ? 8'h37 : _GEN_661; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_663 = 8'h97 == io_in_2 ? 8'h35 : _GEN_662; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_664 = 8'h98 == io_in_2 ? 8'h2b : _GEN_663; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_665 = 8'h99 == io_in_2 ? 8'h29 : _GEN_664; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_666 = 8'h9a == io_in_2 ? 8'h2f : _GEN_665; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_667 = 8'h9b == io_in_2 ? 8'h2d : _GEN_666; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_668 = 8'h9c == io_in_2 ? 8'h23 : _GEN_667; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_669 = 8'h9d == io_in_2 ? 8'h21 : _GEN_668; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_670 = 8'h9e == io_in_2 ? 8'h27 : _GEN_669; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_671 = 8'h9f == io_in_2 ? 8'h25 : _GEN_670; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_672 = 8'ha0 == io_in_2 ? 8'h5b : _GEN_671; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_673 = 8'ha1 == io_in_2 ? 8'h59 : _GEN_672; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_674 = 8'ha2 == io_in_2 ? 8'h5f : _GEN_673; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_675 = 8'ha3 == io_in_2 ? 8'h5d : _GEN_674; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_676 = 8'ha4 == io_in_2 ? 8'h53 : _GEN_675; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_677 = 8'ha5 == io_in_2 ? 8'h51 : _GEN_676; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_678 = 8'ha6 == io_in_2 ? 8'h57 : _GEN_677; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_679 = 8'ha7 == io_in_2 ? 8'h55 : _GEN_678; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_680 = 8'ha8 == io_in_2 ? 8'h4b : _GEN_679; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_681 = 8'ha9 == io_in_2 ? 8'h49 : _GEN_680; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_682 = 8'haa == io_in_2 ? 8'h4f : _GEN_681; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_683 = 8'hab == io_in_2 ? 8'h4d : _GEN_682; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_684 = 8'hac == io_in_2 ? 8'h43 : _GEN_683; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_685 = 8'had == io_in_2 ? 8'h41 : _GEN_684; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_686 = 8'hae == io_in_2 ? 8'h47 : _GEN_685; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_687 = 8'haf == io_in_2 ? 8'h45 : _GEN_686; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_688 = 8'hb0 == io_in_2 ? 8'h7b : _GEN_687; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_689 = 8'hb1 == io_in_2 ? 8'h79 : _GEN_688; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_690 = 8'hb2 == io_in_2 ? 8'h7f : _GEN_689; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_691 = 8'hb3 == io_in_2 ? 8'h7d : _GEN_690; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_692 = 8'hb4 == io_in_2 ? 8'h73 : _GEN_691; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_693 = 8'hb5 == io_in_2 ? 8'h71 : _GEN_692; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_694 = 8'hb6 == io_in_2 ? 8'h77 : _GEN_693; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_695 = 8'hb7 == io_in_2 ? 8'h75 : _GEN_694; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_696 = 8'hb8 == io_in_2 ? 8'h6b : _GEN_695; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_697 = 8'hb9 == io_in_2 ? 8'h69 : _GEN_696; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_698 = 8'hba == io_in_2 ? 8'h6f : _GEN_697; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_699 = 8'hbb == io_in_2 ? 8'h6d : _GEN_698; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_700 = 8'hbc == io_in_2 ? 8'h63 : _GEN_699; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_701 = 8'hbd == io_in_2 ? 8'h61 : _GEN_700; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_702 = 8'hbe == io_in_2 ? 8'h67 : _GEN_701; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_703 = 8'hbf == io_in_2 ? 8'h65 : _GEN_702; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_704 = 8'hc0 == io_in_2 ? 8'h9b : _GEN_703; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_705 = 8'hc1 == io_in_2 ? 8'h99 : _GEN_704; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_706 = 8'hc2 == io_in_2 ? 8'h9f : _GEN_705; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_707 = 8'hc3 == io_in_2 ? 8'h9d : _GEN_706; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_708 = 8'hc4 == io_in_2 ? 8'h93 : _GEN_707; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_709 = 8'hc5 == io_in_2 ? 8'h91 : _GEN_708; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_710 = 8'hc6 == io_in_2 ? 8'h97 : _GEN_709; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_711 = 8'hc7 == io_in_2 ? 8'h95 : _GEN_710; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_712 = 8'hc8 == io_in_2 ? 8'h8b : _GEN_711; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_713 = 8'hc9 == io_in_2 ? 8'h89 : _GEN_712; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_714 = 8'hca == io_in_2 ? 8'h8f : _GEN_713; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_715 = 8'hcb == io_in_2 ? 8'h8d : _GEN_714; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_716 = 8'hcc == io_in_2 ? 8'h83 : _GEN_715; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_717 = 8'hcd == io_in_2 ? 8'h81 : _GEN_716; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_718 = 8'hce == io_in_2 ? 8'h87 : _GEN_717; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_719 = 8'hcf == io_in_2 ? 8'h85 : _GEN_718; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_720 = 8'hd0 == io_in_2 ? 8'hbb : _GEN_719; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_721 = 8'hd1 == io_in_2 ? 8'hb9 : _GEN_720; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_722 = 8'hd2 == io_in_2 ? 8'hbf : _GEN_721; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_723 = 8'hd3 == io_in_2 ? 8'hbd : _GEN_722; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_724 = 8'hd4 == io_in_2 ? 8'hb3 : _GEN_723; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_725 = 8'hd5 == io_in_2 ? 8'hb1 : _GEN_724; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_726 = 8'hd6 == io_in_2 ? 8'hb7 : _GEN_725; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_727 = 8'hd7 == io_in_2 ? 8'hb5 : _GEN_726; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_728 = 8'hd8 == io_in_2 ? 8'hab : _GEN_727; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_729 = 8'hd9 == io_in_2 ? 8'ha9 : _GEN_728; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_730 = 8'hda == io_in_2 ? 8'haf : _GEN_729; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_731 = 8'hdb == io_in_2 ? 8'had : _GEN_730; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_732 = 8'hdc == io_in_2 ? 8'ha3 : _GEN_731; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_733 = 8'hdd == io_in_2 ? 8'ha1 : _GEN_732; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_734 = 8'hde == io_in_2 ? 8'ha7 : _GEN_733; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_735 = 8'hdf == io_in_2 ? 8'ha5 : _GEN_734; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_736 = 8'he0 == io_in_2 ? 8'hdb : _GEN_735; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_737 = 8'he1 == io_in_2 ? 8'hd9 : _GEN_736; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_738 = 8'he2 == io_in_2 ? 8'hdf : _GEN_737; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_739 = 8'he3 == io_in_2 ? 8'hdd : _GEN_738; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_740 = 8'he4 == io_in_2 ? 8'hd3 : _GEN_739; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_741 = 8'he5 == io_in_2 ? 8'hd1 : _GEN_740; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_742 = 8'he6 == io_in_2 ? 8'hd7 : _GEN_741; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_743 = 8'he7 == io_in_2 ? 8'hd5 : _GEN_742; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_744 = 8'he8 == io_in_2 ? 8'hcb : _GEN_743; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_745 = 8'he9 == io_in_2 ? 8'hc9 : _GEN_744; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_746 = 8'hea == io_in_2 ? 8'hcf : _GEN_745; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_747 = 8'heb == io_in_2 ? 8'hcd : _GEN_746; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_748 = 8'hec == io_in_2 ? 8'hc3 : _GEN_747; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_749 = 8'hed == io_in_2 ? 8'hc1 : _GEN_748; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_750 = 8'hee == io_in_2 ? 8'hc7 : _GEN_749; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_751 = 8'hef == io_in_2 ? 8'hc5 : _GEN_750; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_752 = 8'hf0 == io_in_2 ? 8'hfb : _GEN_751; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_753 = 8'hf1 == io_in_2 ? 8'hf9 : _GEN_752; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_754 = 8'hf2 == io_in_2 ? 8'hff : _GEN_753; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_755 = 8'hf3 == io_in_2 ? 8'hfd : _GEN_754; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_756 = 8'hf4 == io_in_2 ? 8'hf3 : _GEN_755; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_757 = 8'hf5 == io_in_2 ? 8'hf1 : _GEN_756; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_758 = 8'hf6 == io_in_2 ? 8'hf7 : _GEN_757; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_759 = 8'hf7 == io_in_2 ? 8'hf5 : _GEN_758; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_760 = 8'hf8 == io_in_2 ? 8'heb : _GEN_759; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_761 = 8'hf9 == io_in_2 ? 8'he9 : _GEN_760; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_762 = 8'hfa == io_in_2 ? 8'hef : _GEN_761; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_763 = 8'hfb == io_in_2 ? 8'hed : _GEN_762; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_764 = 8'hfc == io_in_2 ? 8'he3 : _GEN_763; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_765 = 8'hfd == io_in_2 ? 8'he1 : _GEN_764; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_766 = 8'hfe == io_in_2 ? 8'he7 : _GEN_765; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _GEN_767 = 8'hff == io_in_2 ? 8'he5 : _GEN_766; // @[AES_EncryptionFSM.scala 297:42 AES_EncryptionFSM.scala 297:42]
  wire [7:0] _T_5 = _T_4 ^ _GEN_767; // @[AES_EncryptionFSM.scala 297:42]
  wire [7:0] _T_6 = _T_5 ^ io_in_2; // @[AES_EncryptionFSM.scala 297:59]
  wire [7:0] _T_8 = io_in_0 ^ io_in_1; // @[AES_EncryptionFSM.scala 298:25]
  wire [7:0] _T_9 = _T_8 ^ _GEN_767; // @[AES_EncryptionFSM.scala 298:36]
  wire [7:0] _GEN_769 = 8'h1 == io_in_3 ? 8'h2 : 8'h0; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_770 = 8'h2 == io_in_3 ? 8'h4 : _GEN_769; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_771 = 8'h3 == io_in_3 ? 8'h6 : _GEN_770; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_772 = 8'h4 == io_in_3 ? 8'h8 : _GEN_771; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_773 = 8'h5 == io_in_3 ? 8'ha : _GEN_772; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_774 = 8'h6 == io_in_3 ? 8'hc : _GEN_773; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_775 = 8'h7 == io_in_3 ? 8'he : _GEN_774; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_776 = 8'h8 == io_in_3 ? 8'h10 : _GEN_775; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_777 = 8'h9 == io_in_3 ? 8'h12 : _GEN_776; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_778 = 8'ha == io_in_3 ? 8'h14 : _GEN_777; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_779 = 8'hb == io_in_3 ? 8'h16 : _GEN_778; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_780 = 8'hc == io_in_3 ? 8'h18 : _GEN_779; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_781 = 8'hd == io_in_3 ? 8'h1a : _GEN_780; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_782 = 8'he == io_in_3 ? 8'h1c : _GEN_781; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_783 = 8'hf == io_in_3 ? 8'h1e : _GEN_782; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_784 = 8'h10 == io_in_3 ? 8'h20 : _GEN_783; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_785 = 8'h11 == io_in_3 ? 8'h22 : _GEN_784; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_786 = 8'h12 == io_in_3 ? 8'h24 : _GEN_785; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_787 = 8'h13 == io_in_3 ? 8'h26 : _GEN_786; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_788 = 8'h14 == io_in_3 ? 8'h28 : _GEN_787; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_789 = 8'h15 == io_in_3 ? 8'h2a : _GEN_788; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_790 = 8'h16 == io_in_3 ? 8'h2c : _GEN_789; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_791 = 8'h17 == io_in_3 ? 8'h2e : _GEN_790; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_792 = 8'h18 == io_in_3 ? 8'h30 : _GEN_791; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_793 = 8'h19 == io_in_3 ? 8'h32 : _GEN_792; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_794 = 8'h1a == io_in_3 ? 8'h34 : _GEN_793; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_795 = 8'h1b == io_in_3 ? 8'h36 : _GEN_794; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_796 = 8'h1c == io_in_3 ? 8'h38 : _GEN_795; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_797 = 8'h1d == io_in_3 ? 8'h3a : _GEN_796; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_798 = 8'h1e == io_in_3 ? 8'h3c : _GEN_797; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_799 = 8'h1f == io_in_3 ? 8'h3e : _GEN_798; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_800 = 8'h20 == io_in_3 ? 8'h40 : _GEN_799; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_801 = 8'h21 == io_in_3 ? 8'h42 : _GEN_800; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_802 = 8'h22 == io_in_3 ? 8'h44 : _GEN_801; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_803 = 8'h23 == io_in_3 ? 8'h46 : _GEN_802; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_804 = 8'h24 == io_in_3 ? 8'h48 : _GEN_803; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_805 = 8'h25 == io_in_3 ? 8'h4a : _GEN_804; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_806 = 8'h26 == io_in_3 ? 8'h4c : _GEN_805; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_807 = 8'h27 == io_in_3 ? 8'h4e : _GEN_806; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_808 = 8'h28 == io_in_3 ? 8'h50 : _GEN_807; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_809 = 8'h29 == io_in_3 ? 8'h52 : _GEN_808; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_810 = 8'h2a == io_in_3 ? 8'h54 : _GEN_809; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_811 = 8'h2b == io_in_3 ? 8'h56 : _GEN_810; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_812 = 8'h2c == io_in_3 ? 8'h58 : _GEN_811; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_813 = 8'h2d == io_in_3 ? 8'h5a : _GEN_812; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_814 = 8'h2e == io_in_3 ? 8'h5c : _GEN_813; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_815 = 8'h2f == io_in_3 ? 8'h5e : _GEN_814; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_816 = 8'h30 == io_in_3 ? 8'h60 : _GEN_815; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_817 = 8'h31 == io_in_3 ? 8'h62 : _GEN_816; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_818 = 8'h32 == io_in_3 ? 8'h64 : _GEN_817; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_819 = 8'h33 == io_in_3 ? 8'h66 : _GEN_818; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_820 = 8'h34 == io_in_3 ? 8'h68 : _GEN_819; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_821 = 8'h35 == io_in_3 ? 8'h6a : _GEN_820; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_822 = 8'h36 == io_in_3 ? 8'h6c : _GEN_821; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_823 = 8'h37 == io_in_3 ? 8'h6e : _GEN_822; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_824 = 8'h38 == io_in_3 ? 8'h70 : _GEN_823; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_825 = 8'h39 == io_in_3 ? 8'h72 : _GEN_824; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_826 = 8'h3a == io_in_3 ? 8'h74 : _GEN_825; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_827 = 8'h3b == io_in_3 ? 8'h76 : _GEN_826; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_828 = 8'h3c == io_in_3 ? 8'h78 : _GEN_827; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_829 = 8'h3d == io_in_3 ? 8'h7a : _GEN_828; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_830 = 8'h3e == io_in_3 ? 8'h7c : _GEN_829; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_831 = 8'h3f == io_in_3 ? 8'h7e : _GEN_830; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_832 = 8'h40 == io_in_3 ? 8'h80 : _GEN_831; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_833 = 8'h41 == io_in_3 ? 8'h82 : _GEN_832; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_834 = 8'h42 == io_in_3 ? 8'h84 : _GEN_833; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_835 = 8'h43 == io_in_3 ? 8'h86 : _GEN_834; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_836 = 8'h44 == io_in_3 ? 8'h88 : _GEN_835; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_837 = 8'h45 == io_in_3 ? 8'h8a : _GEN_836; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_838 = 8'h46 == io_in_3 ? 8'h8c : _GEN_837; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_839 = 8'h47 == io_in_3 ? 8'h8e : _GEN_838; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_840 = 8'h48 == io_in_3 ? 8'h90 : _GEN_839; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_841 = 8'h49 == io_in_3 ? 8'h92 : _GEN_840; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_842 = 8'h4a == io_in_3 ? 8'h94 : _GEN_841; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_843 = 8'h4b == io_in_3 ? 8'h96 : _GEN_842; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_844 = 8'h4c == io_in_3 ? 8'h98 : _GEN_843; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_845 = 8'h4d == io_in_3 ? 8'h9a : _GEN_844; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_846 = 8'h4e == io_in_3 ? 8'h9c : _GEN_845; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_847 = 8'h4f == io_in_3 ? 8'h9e : _GEN_846; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_848 = 8'h50 == io_in_3 ? 8'ha0 : _GEN_847; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_849 = 8'h51 == io_in_3 ? 8'ha2 : _GEN_848; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_850 = 8'h52 == io_in_3 ? 8'ha4 : _GEN_849; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_851 = 8'h53 == io_in_3 ? 8'ha6 : _GEN_850; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_852 = 8'h54 == io_in_3 ? 8'ha8 : _GEN_851; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_853 = 8'h55 == io_in_3 ? 8'haa : _GEN_852; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_854 = 8'h56 == io_in_3 ? 8'hac : _GEN_853; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_855 = 8'h57 == io_in_3 ? 8'hae : _GEN_854; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_856 = 8'h58 == io_in_3 ? 8'hb0 : _GEN_855; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_857 = 8'h59 == io_in_3 ? 8'hb2 : _GEN_856; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_858 = 8'h5a == io_in_3 ? 8'hb4 : _GEN_857; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_859 = 8'h5b == io_in_3 ? 8'hb6 : _GEN_858; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_860 = 8'h5c == io_in_3 ? 8'hb8 : _GEN_859; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_861 = 8'h5d == io_in_3 ? 8'hba : _GEN_860; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_862 = 8'h5e == io_in_3 ? 8'hbc : _GEN_861; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_863 = 8'h5f == io_in_3 ? 8'hbe : _GEN_862; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_864 = 8'h60 == io_in_3 ? 8'hc0 : _GEN_863; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_865 = 8'h61 == io_in_3 ? 8'hc2 : _GEN_864; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_866 = 8'h62 == io_in_3 ? 8'hc4 : _GEN_865; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_867 = 8'h63 == io_in_3 ? 8'hc6 : _GEN_866; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_868 = 8'h64 == io_in_3 ? 8'hc8 : _GEN_867; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_869 = 8'h65 == io_in_3 ? 8'hca : _GEN_868; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_870 = 8'h66 == io_in_3 ? 8'hcc : _GEN_869; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_871 = 8'h67 == io_in_3 ? 8'hce : _GEN_870; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_872 = 8'h68 == io_in_3 ? 8'hd0 : _GEN_871; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_873 = 8'h69 == io_in_3 ? 8'hd2 : _GEN_872; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_874 = 8'h6a == io_in_3 ? 8'hd4 : _GEN_873; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_875 = 8'h6b == io_in_3 ? 8'hd6 : _GEN_874; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_876 = 8'h6c == io_in_3 ? 8'hd8 : _GEN_875; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_877 = 8'h6d == io_in_3 ? 8'hda : _GEN_876; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_878 = 8'h6e == io_in_3 ? 8'hdc : _GEN_877; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_879 = 8'h6f == io_in_3 ? 8'hde : _GEN_878; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_880 = 8'h70 == io_in_3 ? 8'he0 : _GEN_879; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_881 = 8'h71 == io_in_3 ? 8'he2 : _GEN_880; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_882 = 8'h72 == io_in_3 ? 8'he4 : _GEN_881; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_883 = 8'h73 == io_in_3 ? 8'he6 : _GEN_882; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_884 = 8'h74 == io_in_3 ? 8'he8 : _GEN_883; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_885 = 8'h75 == io_in_3 ? 8'hea : _GEN_884; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_886 = 8'h76 == io_in_3 ? 8'hec : _GEN_885; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_887 = 8'h77 == io_in_3 ? 8'hee : _GEN_886; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_888 = 8'h78 == io_in_3 ? 8'hf0 : _GEN_887; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_889 = 8'h79 == io_in_3 ? 8'hf2 : _GEN_888; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_890 = 8'h7a == io_in_3 ? 8'hf4 : _GEN_889; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_891 = 8'h7b == io_in_3 ? 8'hf6 : _GEN_890; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_892 = 8'h7c == io_in_3 ? 8'hf8 : _GEN_891; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_893 = 8'h7d == io_in_3 ? 8'hfa : _GEN_892; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_894 = 8'h7e == io_in_3 ? 8'hfc : _GEN_893; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_895 = 8'h7f == io_in_3 ? 8'hfe : _GEN_894; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_896 = 8'h80 == io_in_3 ? 8'h1b : _GEN_895; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_897 = 8'h81 == io_in_3 ? 8'h19 : _GEN_896; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_898 = 8'h82 == io_in_3 ? 8'h1f : _GEN_897; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_899 = 8'h83 == io_in_3 ? 8'h1d : _GEN_898; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_900 = 8'h84 == io_in_3 ? 8'h13 : _GEN_899; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_901 = 8'h85 == io_in_3 ? 8'h11 : _GEN_900; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_902 = 8'h86 == io_in_3 ? 8'h17 : _GEN_901; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_903 = 8'h87 == io_in_3 ? 8'h15 : _GEN_902; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_904 = 8'h88 == io_in_3 ? 8'hb : _GEN_903; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_905 = 8'h89 == io_in_3 ? 8'h9 : _GEN_904; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_906 = 8'h8a == io_in_3 ? 8'hf : _GEN_905; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_907 = 8'h8b == io_in_3 ? 8'hd : _GEN_906; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_908 = 8'h8c == io_in_3 ? 8'h3 : _GEN_907; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_909 = 8'h8d == io_in_3 ? 8'h1 : _GEN_908; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_910 = 8'h8e == io_in_3 ? 8'h7 : _GEN_909; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_911 = 8'h8f == io_in_3 ? 8'h5 : _GEN_910; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_912 = 8'h90 == io_in_3 ? 8'h3b : _GEN_911; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_913 = 8'h91 == io_in_3 ? 8'h39 : _GEN_912; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_914 = 8'h92 == io_in_3 ? 8'h3f : _GEN_913; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_915 = 8'h93 == io_in_3 ? 8'h3d : _GEN_914; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_916 = 8'h94 == io_in_3 ? 8'h33 : _GEN_915; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_917 = 8'h95 == io_in_3 ? 8'h31 : _GEN_916; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_918 = 8'h96 == io_in_3 ? 8'h37 : _GEN_917; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_919 = 8'h97 == io_in_3 ? 8'h35 : _GEN_918; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_920 = 8'h98 == io_in_3 ? 8'h2b : _GEN_919; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_921 = 8'h99 == io_in_3 ? 8'h29 : _GEN_920; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_922 = 8'h9a == io_in_3 ? 8'h2f : _GEN_921; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_923 = 8'h9b == io_in_3 ? 8'h2d : _GEN_922; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_924 = 8'h9c == io_in_3 ? 8'h23 : _GEN_923; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_925 = 8'h9d == io_in_3 ? 8'h21 : _GEN_924; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_926 = 8'h9e == io_in_3 ? 8'h27 : _GEN_925; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_927 = 8'h9f == io_in_3 ? 8'h25 : _GEN_926; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_928 = 8'ha0 == io_in_3 ? 8'h5b : _GEN_927; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_929 = 8'ha1 == io_in_3 ? 8'h59 : _GEN_928; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_930 = 8'ha2 == io_in_3 ? 8'h5f : _GEN_929; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_931 = 8'ha3 == io_in_3 ? 8'h5d : _GEN_930; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_932 = 8'ha4 == io_in_3 ? 8'h53 : _GEN_931; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_933 = 8'ha5 == io_in_3 ? 8'h51 : _GEN_932; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_934 = 8'ha6 == io_in_3 ? 8'h57 : _GEN_933; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_935 = 8'ha7 == io_in_3 ? 8'h55 : _GEN_934; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_936 = 8'ha8 == io_in_3 ? 8'h4b : _GEN_935; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_937 = 8'ha9 == io_in_3 ? 8'h49 : _GEN_936; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_938 = 8'haa == io_in_3 ? 8'h4f : _GEN_937; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_939 = 8'hab == io_in_3 ? 8'h4d : _GEN_938; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_940 = 8'hac == io_in_3 ? 8'h43 : _GEN_939; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_941 = 8'had == io_in_3 ? 8'h41 : _GEN_940; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_942 = 8'hae == io_in_3 ? 8'h47 : _GEN_941; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_943 = 8'haf == io_in_3 ? 8'h45 : _GEN_942; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_944 = 8'hb0 == io_in_3 ? 8'h7b : _GEN_943; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_945 = 8'hb1 == io_in_3 ? 8'h79 : _GEN_944; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_946 = 8'hb2 == io_in_3 ? 8'h7f : _GEN_945; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_947 = 8'hb3 == io_in_3 ? 8'h7d : _GEN_946; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_948 = 8'hb4 == io_in_3 ? 8'h73 : _GEN_947; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_949 = 8'hb5 == io_in_3 ? 8'h71 : _GEN_948; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_950 = 8'hb6 == io_in_3 ? 8'h77 : _GEN_949; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_951 = 8'hb7 == io_in_3 ? 8'h75 : _GEN_950; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_952 = 8'hb8 == io_in_3 ? 8'h6b : _GEN_951; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_953 = 8'hb9 == io_in_3 ? 8'h69 : _GEN_952; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_954 = 8'hba == io_in_3 ? 8'h6f : _GEN_953; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_955 = 8'hbb == io_in_3 ? 8'h6d : _GEN_954; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_956 = 8'hbc == io_in_3 ? 8'h63 : _GEN_955; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_957 = 8'hbd == io_in_3 ? 8'h61 : _GEN_956; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_958 = 8'hbe == io_in_3 ? 8'h67 : _GEN_957; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_959 = 8'hbf == io_in_3 ? 8'h65 : _GEN_958; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_960 = 8'hc0 == io_in_3 ? 8'h9b : _GEN_959; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_961 = 8'hc1 == io_in_3 ? 8'h99 : _GEN_960; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_962 = 8'hc2 == io_in_3 ? 8'h9f : _GEN_961; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_963 = 8'hc3 == io_in_3 ? 8'h9d : _GEN_962; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_964 = 8'hc4 == io_in_3 ? 8'h93 : _GEN_963; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_965 = 8'hc5 == io_in_3 ? 8'h91 : _GEN_964; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_966 = 8'hc6 == io_in_3 ? 8'h97 : _GEN_965; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_967 = 8'hc7 == io_in_3 ? 8'h95 : _GEN_966; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_968 = 8'hc8 == io_in_3 ? 8'h8b : _GEN_967; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_969 = 8'hc9 == io_in_3 ? 8'h89 : _GEN_968; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_970 = 8'hca == io_in_3 ? 8'h8f : _GEN_969; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_971 = 8'hcb == io_in_3 ? 8'h8d : _GEN_970; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_972 = 8'hcc == io_in_3 ? 8'h83 : _GEN_971; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_973 = 8'hcd == io_in_3 ? 8'h81 : _GEN_972; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_974 = 8'hce == io_in_3 ? 8'h87 : _GEN_973; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_975 = 8'hcf == io_in_3 ? 8'h85 : _GEN_974; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_976 = 8'hd0 == io_in_3 ? 8'hbb : _GEN_975; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_977 = 8'hd1 == io_in_3 ? 8'hb9 : _GEN_976; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_978 = 8'hd2 == io_in_3 ? 8'hbf : _GEN_977; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_979 = 8'hd3 == io_in_3 ? 8'hbd : _GEN_978; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_980 = 8'hd4 == io_in_3 ? 8'hb3 : _GEN_979; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_981 = 8'hd5 == io_in_3 ? 8'hb1 : _GEN_980; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_982 = 8'hd6 == io_in_3 ? 8'hb7 : _GEN_981; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_983 = 8'hd7 == io_in_3 ? 8'hb5 : _GEN_982; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_984 = 8'hd8 == io_in_3 ? 8'hab : _GEN_983; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_985 = 8'hd9 == io_in_3 ? 8'ha9 : _GEN_984; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_986 = 8'hda == io_in_3 ? 8'haf : _GEN_985; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_987 = 8'hdb == io_in_3 ? 8'had : _GEN_986; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_988 = 8'hdc == io_in_3 ? 8'ha3 : _GEN_987; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_989 = 8'hdd == io_in_3 ? 8'ha1 : _GEN_988; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_990 = 8'hde == io_in_3 ? 8'ha7 : _GEN_989; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_991 = 8'hdf == io_in_3 ? 8'ha5 : _GEN_990; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_992 = 8'he0 == io_in_3 ? 8'hdb : _GEN_991; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_993 = 8'he1 == io_in_3 ? 8'hd9 : _GEN_992; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_994 = 8'he2 == io_in_3 ? 8'hdf : _GEN_993; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_995 = 8'he3 == io_in_3 ? 8'hdd : _GEN_994; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_996 = 8'he4 == io_in_3 ? 8'hd3 : _GEN_995; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_997 = 8'he5 == io_in_3 ? 8'hd1 : _GEN_996; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_998 = 8'he6 == io_in_3 ? 8'hd7 : _GEN_997; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_999 = 8'he7 == io_in_3 ? 8'hd5 : _GEN_998; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1000 = 8'he8 == io_in_3 ? 8'hcb : _GEN_999; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1001 = 8'he9 == io_in_3 ? 8'hc9 : _GEN_1000; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1002 = 8'hea == io_in_3 ? 8'hcf : _GEN_1001; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1003 = 8'heb == io_in_3 ? 8'hcd : _GEN_1002; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1004 = 8'hec == io_in_3 ? 8'hc3 : _GEN_1003; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1005 = 8'hed == io_in_3 ? 8'hc1 : _GEN_1004; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1006 = 8'hee == io_in_3 ? 8'hc7 : _GEN_1005; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1007 = 8'hef == io_in_3 ? 8'hc5 : _GEN_1006; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1008 = 8'hf0 == io_in_3 ? 8'hfb : _GEN_1007; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1009 = 8'hf1 == io_in_3 ? 8'hf9 : _GEN_1008; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1010 = 8'hf2 == io_in_3 ? 8'hff : _GEN_1009; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1011 = 8'hf3 == io_in_3 ? 8'hfd : _GEN_1010; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1012 = 8'hf4 == io_in_3 ? 8'hf3 : _GEN_1011; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1013 = 8'hf5 == io_in_3 ? 8'hf1 : _GEN_1012; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1014 = 8'hf6 == io_in_3 ? 8'hf7 : _GEN_1013; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1015 = 8'hf7 == io_in_3 ? 8'hf5 : _GEN_1014; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1016 = 8'hf8 == io_in_3 ? 8'heb : _GEN_1015; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1017 = 8'hf9 == io_in_3 ? 8'he9 : _GEN_1016; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1018 = 8'hfa == io_in_3 ? 8'hef : _GEN_1017; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1019 = 8'hfb == io_in_3 ? 8'hed : _GEN_1018; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1020 = 8'hfc == io_in_3 ? 8'he3 : _GEN_1019; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1021 = 8'hfd == io_in_3 ? 8'he1 : _GEN_1020; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1022 = 8'hfe == io_in_3 ? 8'he7 : _GEN_1021; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _GEN_1023 = 8'hff == io_in_3 ? 8'he5 : _GEN_1022; // @[AES_EncryptionFSM.scala 298:53 AES_EncryptionFSM.scala 298:53]
  wire [7:0] _T_10 = _T_9 ^ _GEN_1023; // @[AES_EncryptionFSM.scala 298:53]
  wire [7:0] _T_12 = _GEN_255 ^ io_in_0; // @[AES_EncryptionFSM.scala 299:31]
  wire [7:0] _T_13 = _T_12 ^ io_in_1; // @[AES_EncryptionFSM.scala 299:42]
  wire [7:0] _T_14 = _T_13 ^ io_in_2; // @[AES_EncryptionFSM.scala 299:53]
  assign io_out_0 = _T_2 ^ io_in_3; // @[AES_EncryptionFSM.scala 296:70]
  assign io_out_1 = _T_6 ^ io_in_3; // @[AES_EncryptionFSM.scala 297:70]
  assign io_out_2 = _T_10 ^ io_in_3; // @[AES_EncryptionFSM.scala 298:70]
  assign io_out_3 = _T_14 ^ _GEN_1023; // @[AES_EncryptionFSM.scala 299:64]
endmodule
module AES_MixColumns(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3
);
  wire [7:0] PEs_0_io_in_0; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_0_io_in_1; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_0_io_in_2; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_0_io_in_3; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_0_io_out_0; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_0_io_out_1; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_0_io_out_2; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_0_io_out_3; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_1_io_in_0; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_1_io_in_1; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_1_io_in_2; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_1_io_in_3; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_1_io_out_0; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_1_io_out_1; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_1_io_out_2; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_1_io_out_3; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_2_io_in_0; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_2_io_in_1; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_2_io_in_2; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_2_io_in_3; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_2_io_out_0; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_2_io_out_1; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_2_io_out_2; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_2_io_out_3; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_3_io_in_0; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_3_io_in_1; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_3_io_in_2; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_3_io_in_3; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_3_io_out_0; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_3_io_out_1; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_3_io_out_2; // @[AES_EncryptionFSM.scala 246:20]
  wire [7:0] PEs_3_io_out_3; // @[AES_EncryptionFSM.scala 246:20]
  AES_MixColumn PEs_0 ( // @[AES_EncryptionFSM.scala 246:20]
    .io_in_0(PEs_0_io_in_0),
    .io_in_1(PEs_0_io_in_1),
    .io_in_2(PEs_0_io_in_2),
    .io_in_3(PEs_0_io_in_3),
    .io_out_0(PEs_0_io_out_0),
    .io_out_1(PEs_0_io_out_1),
    .io_out_2(PEs_0_io_out_2),
    .io_out_3(PEs_0_io_out_3)
  );
  AES_MixColumn PEs_1 ( // @[AES_EncryptionFSM.scala 246:20]
    .io_in_0(PEs_1_io_in_0),
    .io_in_1(PEs_1_io_in_1),
    .io_in_2(PEs_1_io_in_2),
    .io_in_3(PEs_1_io_in_3),
    .io_out_0(PEs_1_io_out_0),
    .io_out_1(PEs_1_io_out_1),
    .io_out_2(PEs_1_io_out_2),
    .io_out_3(PEs_1_io_out_3)
  );
  AES_MixColumn PEs_2 ( // @[AES_EncryptionFSM.scala 246:20]
    .io_in_0(PEs_2_io_in_0),
    .io_in_1(PEs_2_io_in_1),
    .io_in_2(PEs_2_io_in_2),
    .io_in_3(PEs_2_io_in_3),
    .io_out_0(PEs_2_io_out_0),
    .io_out_1(PEs_2_io_out_1),
    .io_out_2(PEs_2_io_out_2),
    .io_out_3(PEs_2_io_out_3)
  );
  AES_MixColumn PEs_3 ( // @[AES_EncryptionFSM.scala 246:20]
    .io_in_0(PEs_3_io_in_0),
    .io_in_1(PEs_3_io_in_1),
    .io_in_2(PEs_3_io_in_2),
    .io_in_3(PEs_3_io_in_3),
    .io_out_0(PEs_3_io_out_0),
    .io_out_1(PEs_3_io_out_1),
    .io_out_2(PEs_3_io_out_2),
    .io_out_3(PEs_3_io_out_3)
  );
  assign io_out_state_0_0 = PEs_0_io_out_0; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_0_1 = PEs_0_io_out_1; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_0_2 = PEs_0_io_out_2; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_0_3 = PEs_0_io_out_3; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_1_0 = PEs_1_io_out_0; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_1_1 = PEs_1_io_out_1; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_1_2 = PEs_1_io_out_2; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_1_3 = PEs_1_io_out_3; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_2_0 = PEs_2_io_out_0; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_2_1 = PEs_2_io_out_1; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_2_2 = PEs_2_io_out_2; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_2_3 = PEs_2_io_out_3; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_3_0 = PEs_3_io_out_0; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_3_1 = PEs_3_io_out_1; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_3_2 = PEs_3_io_out_2; // @[AES_EncryptionFSM.scala 253:21]
  assign io_out_state_3_3 = PEs_3_io_out_3; // @[AES_EncryptionFSM.scala 253:21]
  assign PEs_0_io_in_0 = io_in_state_0_0; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_0_io_in_1 = io_in_state_0_1; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_0_io_in_2 = io_in_state_0_2; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_0_io_in_3 = io_in_state_0_3; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_1_io_in_0 = io_in_state_1_0; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_1_io_in_1 = io_in_state_1_1; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_1_io_in_2 = io_in_state_1_2; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_1_io_in_3 = io_in_state_1_3; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_2_io_in_0 = io_in_state_2_0; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_2_io_in_1 = io_in_state_2_1; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_2_io_in_2 = io_in_state_2_2; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_2_io_in_3 = io_in_state_2_3; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_3_io_in_0 = io_in_state_3_0; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_3_io_in_1 = io_in_state_3_1; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_3_io_in_2 = io_in_state_3_2; // @[AES_EncryptionFSM.scala 252:18]
  assign PEs_3_io_in_3 = io_in_state_3_3; // @[AES_EncryptionFSM.scala 252:18]
endmodule
module AES_RotWord(
  output [31:0] io_out,
  input  [31:0] io_in
);
  wire [23:0] hi = io_in[23:0]; // @[AES_EncryptionFSM.scala 234:22]
  wire [7:0] lo = io_in[31:24]; // @[AES_EncryptionFSM.scala 234:35]
  assign io_out = {hi,lo}; // @[Cat.scala 30:58]
endmodule
module AES_SubWord(
  output [31:0] io_out,
  input  [31:0] io_in
);
  wire [7:0] PEs_0_io_in; // @[AES_EncryptionFSM.scala 220:20]
  wire [7:0] PEs_0_io_out; // @[AES_EncryptionFSM.scala 220:20]
  wire [7:0] PEs_1_io_in; // @[AES_EncryptionFSM.scala 220:20]
  wire [7:0] PEs_1_io_out; // @[AES_EncryptionFSM.scala 220:20]
  wire [7:0] PEs_2_io_in; // @[AES_EncryptionFSM.scala 220:20]
  wire [7:0] PEs_2_io_out; // @[AES_EncryptionFSM.scala 220:20]
  wire [7:0] PEs_3_io_in; // @[AES_EncryptionFSM.scala 220:20]
  wire [7:0] PEs_3_io_out; // @[AES_EncryptionFSM.scala 220:20]
  wire [15:0] lo = {PEs_1_io_out,PEs_0_io_out}; // @[Cat.scala 30:58]
  wire [15:0] hi = {PEs_3_io_out,PEs_2_io_out}; // @[Cat.scala 30:58]
  AES_S PEs_0 ( // @[AES_EncryptionFSM.scala 220:20]
    .io_in(PEs_0_io_in),
    .io_out(PEs_0_io_out)
  );
  AES_S PEs_1 ( // @[AES_EncryptionFSM.scala 220:20]
    .io_in(PEs_1_io_in),
    .io_out(PEs_1_io_out)
  );
  AES_S PEs_2 ( // @[AES_EncryptionFSM.scala 220:20]
    .io_in(PEs_2_io_in),
    .io_out(PEs_2_io_out)
  );
  AES_S PEs_3 ( // @[AES_EncryptionFSM.scala 220:20]
    .io_in(PEs_3_io_in),
    .io_out(PEs_3_io_out)
  );
  assign io_out = {hi,lo}; // @[Cat.scala 30:58]
  assign PEs_0_io_in = io_in[7:0]; // @[AES_EncryptionFSM.scala 221:22]
  assign PEs_1_io_in = io_in[15:8]; // @[AES_EncryptionFSM.scala 221:22]
  assign PEs_2_io_in = io_in[23:16]; // @[AES_EncryptionFSM.scala 221:22]
  assign PEs_3_io_in = io_in[31:24]; // @[AES_EncryptionFSM.scala 221:22]
endmodule
module AES_GetNewKey(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3,
  input  [3:0] io_round
);
  wire [31:0] rot_io_out; // @[AES_EncryptionFSM.scala 158:19]
  wire [31:0] rot_io_in; // @[AES_EncryptionFSM.scala 158:19]
  wire [31:0] sub_io_out; // @[AES_EncryptionFSM.scala 161:19]
  wire [31:0] sub_io_in; // @[AES_EncryptionFSM.scala 161:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire  _T_4 = 4'h0 == io_round; // @[Conditional.scala 37:30]
  wire  _T_5 = 4'h1 == io_round; // @[Conditional.scala 37:30]
  wire  _T_6 = 4'h2 == io_round; // @[Conditional.scala 37:30]
  wire  _T_7 = 4'h3 == io_round; // @[Conditional.scala 37:30]
  wire  _T_8 = 4'h4 == io_round; // @[Conditional.scala 37:30]
  wire  _T_9 = 4'h5 == io_round; // @[Conditional.scala 37:30]
  wire  _T_10 = 4'h6 == io_round; // @[Conditional.scala 37:30]
  wire  _T_11 = 4'h7 == io_round; // @[Conditional.scala 37:30]
  wire  _T_12 = 4'h8 == io_round; // @[Conditional.scala 37:30]
  wire  _T_13 = 4'h9 == io_round; // @[Conditional.scala 37:30]
  wire [29:0] _GEN_0 = _T_13 ? 30'h36000000 : 30'h0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 195:12 AES_EncryptionFSM.scala 165:8]
  wire [29:0] _GEN_1 = _T_12 ? 30'h1b000000 : _GEN_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 192:12]
  wire [31:0] _GEN_2 = _T_11 ? 32'h80000000 : {{2'd0}, _GEN_1}; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 189:12]
  wire [31:0] _GEN_3 = _T_10 ? 32'h40000000 : _GEN_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 186:12]
  wire [31:0] _GEN_4 = _T_9 ? 32'h20000000 : _GEN_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 183:12]
  wire [31:0] _GEN_5 = _T_8 ? 32'h10000000 : _GEN_4; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 180:12]
  wire [31:0] _GEN_6 = _T_7 ? 32'h8000000 : _GEN_5; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 177:12]
  wire [31:0] _GEN_7 = _T_6 ? 32'h4000000 : _GEN_6; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 174:12]
  wire [31:0] _GEN_8 = _T_5 ? 32'h2000000 : _GEN_7; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 171:12]
  wire [31:0] Rcon = _T_4 ? 32'h1000000 : _GEN_8; // @[Conditional.scala 40:58 AES_EncryptionFSM.scala 168:12]
  wire [31:0] _T_14 = sub_io_out ^ Rcon; // @[AES_EncryptionFSM.scala 200:20]
  wire [31:0] w5 = _T_14 ^ w0; // @[AES_EncryptionFSM.scala 200:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_EncryptionFSM.scala 201:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_EncryptionFSM.scala 202:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_EncryptionFSM.scala 203:12]
  AES_RotWord rot ( // @[AES_EncryptionFSM.scala 158:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_EncryptionFSM.scala 161:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_EncryptionFSM.scala 206:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_EncryptionFSM.scala 206:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_EncryptionFSM.scala 206:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_EncryptionFSM.scala 206:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_EncryptionFSM.scala 207:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_EncryptionFSM.scala 207:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_EncryptionFSM.scala 207:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_EncryptionFSM.scala 207:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_EncryptionFSM.scala 208:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_EncryptionFSM.scala 208:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_EncryptionFSM.scala 208:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_EncryptionFSM.scala 208:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_EncryptionFSM.scala 209:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_EncryptionFSM.scala 209:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_EncryptionFSM.scala 209:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_EncryptionFSM.scala 209:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_EncryptionFSM.scala 162:13]
endmodule
module AES_ProcessingElement(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3,
  input  [3:0] io_round
);
  wire [7:0] sub_io_out_state_0_0; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_EncryptionFSM.scala 116:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_EncryptionFSM.scala 124:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_EncryptionFSM.scala 127:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_EncryptionFSM.scala 136:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_EncryptionFSM.scala 136:19]
  wire [3:0] key_io_round; // @[AES_EncryptionFSM.scala 136:19]
  AES_SubBytes sub ( // @[AES_EncryptionFSM.scala 116:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_EncryptionFSM.scala 124:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_EncryptionFSM.scala 127:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey key ( // @[AES_EncryptionFSM.scala 136:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3),
    .io_round(key_io_round)
  );
  assign io_out_state_0_0 = io_round == 4'h9 ? shift_io_out_state_0_0 : mix_io_out_state_0_0; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_0_1 = io_round == 4'h9 ? shift_io_out_state_0_1 : mix_io_out_state_0_1; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_0_2 = io_round == 4'h9 ? shift_io_out_state_0_2 : mix_io_out_state_0_2; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_0_3 = io_round == 4'h9 ? shift_io_out_state_0_3 : mix_io_out_state_0_3; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_1_0 = io_round == 4'h9 ? shift_io_out_state_1_0 : mix_io_out_state_1_0; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_1_1 = io_round == 4'h9 ? shift_io_out_state_1_1 : mix_io_out_state_1_1; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_1_2 = io_round == 4'h9 ? shift_io_out_state_1_2 : mix_io_out_state_1_2; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_1_3 = io_round == 4'h9 ? shift_io_out_state_1_3 : mix_io_out_state_1_3; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_2_0 = io_round == 4'h9 ? shift_io_out_state_2_0 : mix_io_out_state_2_0; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_2_1 = io_round == 4'h9 ? shift_io_out_state_2_1 : mix_io_out_state_2_1; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_2_2 = io_round == 4'h9 ? shift_io_out_state_2_2 : mix_io_out_state_2_2; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_2_3 = io_round == 4'h9 ? shift_io_out_state_2_3 : mix_io_out_state_2_3; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_3_0 = io_round == 4'h9 ? shift_io_out_state_3_0 : mix_io_out_state_3_0; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_3_1 = io_round == 4'h9 ? shift_io_out_state_3_1 : mix_io_out_state_3_1; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_3_2 = io_round == 4'h9 ? shift_io_out_state_3_2 : mix_io_out_state_3_2; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_state_3_3 = io_round == 4'h9 ? shift_io_out_state_3_3 : mix_io_out_state_3_3; // @[AES_EncryptionFSM.scala 130:26 AES_EncryptionFSM.scala 131:18 AES_EncryptionFSM.scala 133:18]
  assign io_out_key_0_0 = key_io_out_key_0_0; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_0_1 = key_io_out_key_0_1; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_0_2 = key_io_out_key_0_2; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_0_3 = key_io_out_key_0_3; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_1_0 = key_io_out_key_1_0; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_1_1 = key_io_out_key_1_1; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_1_2 = key_io_out_key_1_2; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_1_3 = key_io_out_key_1_3; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_2_0 = key_io_out_key_2_0; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_2_1 = key_io_out_key_2_1; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_2_2 = key_io_out_key_2_2; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_2_3 = key_io_out_key_2_3; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_3_0 = key_io_out_key_3_0; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_3_1 = key_io_out_key_3_1; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_3_2 = key_io_out_key_3_2; // @[AES_EncryptionFSM.scala 140:14]
  assign io_out_key_3_3 = key_io_out_key_3_3; // @[AES_EncryptionFSM.scala 140:14]
  assign sub_io_in_state_0_0 = io_in_state_0_0 ^ io_in_key_0_0; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_0_1 = io_in_state_0_1 ^ io_in_key_0_1; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_0_2 = io_in_state_0_2 ^ io_in_key_0_2; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_0_3 = io_in_state_0_3 ^ io_in_key_0_3; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_1_0 = io_in_state_1_0 ^ io_in_key_1_0; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_1_1 = io_in_state_1_1 ^ io_in_key_1_1; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_1_2 = io_in_state_1_2 ^ io_in_key_1_2; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_1_3 = io_in_state_1_3 ^ io_in_key_1_3; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_2_0 = io_in_state_2_0 ^ io_in_key_2_0; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_2_1 = io_in_state_2_1 ^ io_in_key_2_1; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_2_2 = io_in_state_2_2 ^ io_in_key_2_2; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_2_3 = io_in_state_2_3 ^ io_in_key_2_3; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_3_0 = io_in_state_3_0 ^ io_in_key_3_0; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_3_1 = io_in_state_3_1 ^ io_in_key_3_1; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_3_2 = io_in_state_3_2 ^ io_in_key_3_2; // @[AES_EncryptionFSM.scala 120:50]
  assign sub_io_in_state_3_3 = io_in_state_3_3 ^ io_in_key_3_3; // @[AES_EncryptionFSM.scala 120:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_EncryptionFSM.scala 125:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_EncryptionFSM.scala 125:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_EncryptionFSM.scala 128:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_EncryptionFSM.scala 128:13]
  assign key_io_in_key_0_0 = io_in_key_0_0; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_0_1 = io_in_key_0_1; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_0_2 = io_in_key_0_2; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_0_3 = io_in_key_0_3; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_1_0 = io_in_key_1_0; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_1_1 = io_in_key_1_1; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_1_2 = io_in_key_1_2; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_1_3 = io_in_key_1_3; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_2_0 = io_in_key_2_0; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_2_1 = io_in_key_2_1; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_2_2 = io_in_key_2_2; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_2_3 = io_in_key_2_3; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_3_0 = io_in_key_3_0; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_3_1 = io_in_key_3_1; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_3_2 = io_in_key_3_2; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_in_key_3_3 = io_in_key_3_3; // @[AES_EncryptionFSM.scala 138:17]
  assign key_io_round = io_round; // @[AES_EncryptionFSM.scala 139:16]
endmodule
module AES_EncryptionFSM(
  input          clock,
  input          reset,
  input          io_out_ready,
  output         io_out_valid,
  output [127:0] io_out_bits_text,
  output [127:0] io_out_bits_key,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits_text,
  input  [127:0] io_in_bits_key
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] initialOp_io_text; // @[AES_EncryptionFSM.scala 24:25]
  wire [127:0] initialOp_io_key; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_0_0; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_0_1; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_0_2; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_0_3; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_1_0; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_1_1; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_1_2; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_1_3; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_2_0; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_2_1; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_2_2; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_2_3; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_3_0; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_3_1; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_3_2; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_state_3_3; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_0_0; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_0_1; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_0_2; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_0_3; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_1_0; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_1_1; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_1_2; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_1_3; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_2_0; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_2_1; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_2_2; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_2_3; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_3_0; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_3_1; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_3_2; // @[AES_EncryptionFSM.scala 24:25]
  wire [7:0] initialOp_io_out_key_3_3; // @[AES_EncryptionFSM.scala 24:25]
  wire [127:0] finalOp_io_out_text; // @[AES_EncryptionFSM.scala 27:23]
  wire [127:0] finalOp_io_out_key; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_0_0; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_0_1; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_0_2; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_0_3; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_1_0; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_1_1; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_1_2; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_1_3; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_2_0; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_2_1; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_2_2; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_2_3; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_3_0; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_3_1; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_3_2; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_state_3_3; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_0_0; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_0_1; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_0_2; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_0_3; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_1_0; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_1_1; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_1_2; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_1_3; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_2_0; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_2_1; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_2_2; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_2_3; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_3_0; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_3_1; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_3_2; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] finalOp_io_in_key_3_3; // @[AES_EncryptionFSM.scala 27:23]
  wire [7:0] pe_io_out_state_0_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_0_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_0_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_0_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_1_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_1_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_1_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_1_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_2_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_2_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_2_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_2_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_3_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_3_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_3_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_state_3_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_0_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_0_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_0_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_0_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_1_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_1_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_1_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_1_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_2_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_2_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_2_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_2_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_3_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_3_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_3_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_out_key_3_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_0_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_0_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_0_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_0_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_1_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_1_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_1_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_1_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_2_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_2_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_2_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_2_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_3_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_3_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_3_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_state_3_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_0_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_0_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_0_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_0_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_1_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_1_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_1_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_1_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_2_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_2_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_2_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_2_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_3_0; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_3_1; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_3_2; // @[AES_EncryptionFSM.scala 30:18]
  wire [7:0] pe_io_in_key_3_3; // @[AES_EncryptionFSM.scala 30:18]
  wire [3:0] pe_io_round; // @[AES_EncryptionFSM.scala 30:18]
  reg [2:0] stateReg; // @[AES_EncryptionFSM.scala 13:25]
  reg [3:0] roundReg; // @[AES_EncryptionFSM.scala 14:25]
  reg [127:0] textReg; // @[AES_EncryptionFSM.scala 15:24]
  reg [127:0] keyReg; // @[AES_EncryptionFSM.scala 16:23]
  reg [7:0] dataReg_state_0_0; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_0_1; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_0_2; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_0_3; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_1_0; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_1_1; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_1_2; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_1_3; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_2_0; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_2_1; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_2_2; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_2_3; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_3_0; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_3_1; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_3_2; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_state_3_3; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_0_0; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_0_1; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_0_2; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_0_3; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_1_0; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_1_1; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_1_2; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_1_3; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_2_0; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_2_1; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_2_2; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_2_3; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_3_0; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_3_1; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_3_2; // @[AES_EncryptionFSM.scala 17:24]
  reg [7:0] dataReg_key_3_3; // @[AES_EncryptionFSM.scala 17:24]
  reg [127:0] resultsReg_text; // @[AES_EncryptionFSM.scala 18:27]
  reg [127:0] resultsReg_key; // @[AES_EncryptionFSM.scala 18:27]
  wire  _T_2 = 3'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h2 == stateReg; // @[Conditional.scala 37:30]
  wire [3:0] _T_6 = roundReg + 4'h1; // @[AES_EncryptionFSM.scala 52:28]
  wire [2:0] _GEN_3 = roundReg == 4'h9 ? 3'h3 : stateReg; // @[AES_EncryptionFSM.scala 53:30 AES_EncryptionFSM.scala 54:18 AES_EncryptionFSM.scala 13:25]
  wire  _T_8 = 3'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h4 == stateReg; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_4 = io_out_ready ? 3'h0 : stateReg; // @[AES_EncryptionFSM.scala 63:26 AES_EncryptionFSM.scala 64:18 AES_EncryptionFSM.scala 13:25]
  wire [2:0] _GEN_5 = _T_9 ? _GEN_4 : stateReg; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 13:25]
  wire [127:0] _GEN_38 = _T_8 ? finalOp_io_out_key : resultsReg_key; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 59:18 AES_EncryptionFSM.scala 18:27]
  wire [127:0] _GEN_39 = _T_8 ? finalOp_io_out_text : resultsReg_text; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 59:18 AES_EncryptionFSM.scala 18:27]
  wire [2:0] _GEN_40 = _T_8 ? 3'h4 : _GEN_5; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 60:16]
  AES_InitialOperation initialOp ( // @[AES_EncryptionFSM.scala 24:25]
    .io_text(initialOp_io_text),
    .io_key(initialOp_io_key),
    .io_out_state_0_0(initialOp_io_out_state_0_0),
    .io_out_state_0_1(initialOp_io_out_state_0_1),
    .io_out_state_0_2(initialOp_io_out_state_0_2),
    .io_out_state_0_3(initialOp_io_out_state_0_3),
    .io_out_state_1_0(initialOp_io_out_state_1_0),
    .io_out_state_1_1(initialOp_io_out_state_1_1),
    .io_out_state_1_2(initialOp_io_out_state_1_2),
    .io_out_state_1_3(initialOp_io_out_state_1_3),
    .io_out_state_2_0(initialOp_io_out_state_2_0),
    .io_out_state_2_1(initialOp_io_out_state_2_1),
    .io_out_state_2_2(initialOp_io_out_state_2_2),
    .io_out_state_2_3(initialOp_io_out_state_2_3),
    .io_out_state_3_0(initialOp_io_out_state_3_0),
    .io_out_state_3_1(initialOp_io_out_state_3_1),
    .io_out_state_3_2(initialOp_io_out_state_3_2),
    .io_out_state_3_3(initialOp_io_out_state_3_3),
    .io_out_key_0_0(initialOp_io_out_key_0_0),
    .io_out_key_0_1(initialOp_io_out_key_0_1),
    .io_out_key_0_2(initialOp_io_out_key_0_2),
    .io_out_key_0_3(initialOp_io_out_key_0_3),
    .io_out_key_1_0(initialOp_io_out_key_1_0),
    .io_out_key_1_1(initialOp_io_out_key_1_1),
    .io_out_key_1_2(initialOp_io_out_key_1_2),
    .io_out_key_1_3(initialOp_io_out_key_1_3),
    .io_out_key_2_0(initialOp_io_out_key_2_0),
    .io_out_key_2_1(initialOp_io_out_key_2_1),
    .io_out_key_2_2(initialOp_io_out_key_2_2),
    .io_out_key_2_3(initialOp_io_out_key_2_3),
    .io_out_key_3_0(initialOp_io_out_key_3_0),
    .io_out_key_3_1(initialOp_io_out_key_3_1),
    .io_out_key_3_2(initialOp_io_out_key_3_2),
    .io_out_key_3_3(initialOp_io_out_key_3_3)
  );
  AES_FinalOperation finalOp ( // @[AES_EncryptionFSM.scala 27:23]
    .io_out_text(finalOp_io_out_text),
    .io_out_key(finalOp_io_out_key),
    .io_in_state_0_0(finalOp_io_in_state_0_0),
    .io_in_state_0_1(finalOp_io_in_state_0_1),
    .io_in_state_0_2(finalOp_io_in_state_0_2),
    .io_in_state_0_3(finalOp_io_in_state_0_3),
    .io_in_state_1_0(finalOp_io_in_state_1_0),
    .io_in_state_1_1(finalOp_io_in_state_1_1),
    .io_in_state_1_2(finalOp_io_in_state_1_2),
    .io_in_state_1_3(finalOp_io_in_state_1_3),
    .io_in_state_2_0(finalOp_io_in_state_2_0),
    .io_in_state_2_1(finalOp_io_in_state_2_1),
    .io_in_state_2_2(finalOp_io_in_state_2_2),
    .io_in_state_2_3(finalOp_io_in_state_2_3),
    .io_in_state_3_0(finalOp_io_in_state_3_0),
    .io_in_state_3_1(finalOp_io_in_state_3_1),
    .io_in_state_3_2(finalOp_io_in_state_3_2),
    .io_in_state_3_3(finalOp_io_in_state_3_3),
    .io_in_key_0_0(finalOp_io_in_key_0_0),
    .io_in_key_0_1(finalOp_io_in_key_0_1),
    .io_in_key_0_2(finalOp_io_in_key_0_2),
    .io_in_key_0_3(finalOp_io_in_key_0_3),
    .io_in_key_1_0(finalOp_io_in_key_1_0),
    .io_in_key_1_1(finalOp_io_in_key_1_1),
    .io_in_key_1_2(finalOp_io_in_key_1_2),
    .io_in_key_1_3(finalOp_io_in_key_1_3),
    .io_in_key_2_0(finalOp_io_in_key_2_0),
    .io_in_key_2_1(finalOp_io_in_key_2_1),
    .io_in_key_2_2(finalOp_io_in_key_2_2),
    .io_in_key_2_3(finalOp_io_in_key_2_3),
    .io_in_key_3_0(finalOp_io_in_key_3_0),
    .io_in_key_3_1(finalOp_io_in_key_3_1),
    .io_in_key_3_2(finalOp_io_in_key_3_2),
    .io_in_key_3_3(finalOp_io_in_key_3_3)
  );
  AES_ProcessingElement pe ( // @[AES_EncryptionFSM.scala 30:18]
    .io_out_state_0_0(pe_io_out_state_0_0),
    .io_out_state_0_1(pe_io_out_state_0_1),
    .io_out_state_0_2(pe_io_out_state_0_2),
    .io_out_state_0_3(pe_io_out_state_0_3),
    .io_out_state_1_0(pe_io_out_state_1_0),
    .io_out_state_1_1(pe_io_out_state_1_1),
    .io_out_state_1_2(pe_io_out_state_1_2),
    .io_out_state_1_3(pe_io_out_state_1_3),
    .io_out_state_2_0(pe_io_out_state_2_0),
    .io_out_state_2_1(pe_io_out_state_2_1),
    .io_out_state_2_2(pe_io_out_state_2_2),
    .io_out_state_2_3(pe_io_out_state_2_3),
    .io_out_state_3_0(pe_io_out_state_3_0),
    .io_out_state_3_1(pe_io_out_state_3_1),
    .io_out_state_3_2(pe_io_out_state_3_2),
    .io_out_state_3_3(pe_io_out_state_3_3),
    .io_out_key_0_0(pe_io_out_key_0_0),
    .io_out_key_0_1(pe_io_out_key_0_1),
    .io_out_key_0_2(pe_io_out_key_0_2),
    .io_out_key_0_3(pe_io_out_key_0_3),
    .io_out_key_1_0(pe_io_out_key_1_0),
    .io_out_key_1_1(pe_io_out_key_1_1),
    .io_out_key_1_2(pe_io_out_key_1_2),
    .io_out_key_1_3(pe_io_out_key_1_3),
    .io_out_key_2_0(pe_io_out_key_2_0),
    .io_out_key_2_1(pe_io_out_key_2_1),
    .io_out_key_2_2(pe_io_out_key_2_2),
    .io_out_key_2_3(pe_io_out_key_2_3),
    .io_out_key_3_0(pe_io_out_key_3_0),
    .io_out_key_3_1(pe_io_out_key_3_1),
    .io_out_key_3_2(pe_io_out_key_3_2),
    .io_out_key_3_3(pe_io_out_key_3_3),
    .io_in_state_0_0(pe_io_in_state_0_0),
    .io_in_state_0_1(pe_io_in_state_0_1),
    .io_in_state_0_2(pe_io_in_state_0_2),
    .io_in_state_0_3(pe_io_in_state_0_3),
    .io_in_state_1_0(pe_io_in_state_1_0),
    .io_in_state_1_1(pe_io_in_state_1_1),
    .io_in_state_1_2(pe_io_in_state_1_2),
    .io_in_state_1_3(pe_io_in_state_1_3),
    .io_in_state_2_0(pe_io_in_state_2_0),
    .io_in_state_2_1(pe_io_in_state_2_1),
    .io_in_state_2_2(pe_io_in_state_2_2),
    .io_in_state_2_3(pe_io_in_state_2_3),
    .io_in_state_3_0(pe_io_in_state_3_0),
    .io_in_state_3_1(pe_io_in_state_3_1),
    .io_in_state_3_2(pe_io_in_state_3_2),
    .io_in_state_3_3(pe_io_in_state_3_3),
    .io_in_key_0_0(pe_io_in_key_0_0),
    .io_in_key_0_1(pe_io_in_key_0_1),
    .io_in_key_0_2(pe_io_in_key_0_2),
    .io_in_key_0_3(pe_io_in_key_0_3),
    .io_in_key_1_0(pe_io_in_key_1_0),
    .io_in_key_1_1(pe_io_in_key_1_1),
    .io_in_key_1_2(pe_io_in_key_1_2),
    .io_in_key_1_3(pe_io_in_key_1_3),
    .io_in_key_2_0(pe_io_in_key_2_0),
    .io_in_key_2_1(pe_io_in_key_2_1),
    .io_in_key_2_2(pe_io_in_key_2_2),
    .io_in_key_2_3(pe_io_in_key_2_3),
    .io_in_key_3_0(pe_io_in_key_3_0),
    .io_in_key_3_1(pe_io_in_key_3_1),
    .io_in_key_3_2(pe_io_in_key_3_2),
    .io_in_key_3_3(pe_io_in_key_3_3),
    .io_round(pe_io_round)
  );
  assign io_out_valid = stateReg == 3'h4; // @[AES_EncryptionFSM.scala 21:28]
  assign io_out_bits_text = resultsReg_text; // @[AES_EncryptionFSM.scala 22:15]
  assign io_out_bits_key = resultsReg_key; // @[AES_EncryptionFSM.scala 22:15]
  assign io_in_ready = stateReg == 3'h0; // @[AES_EncryptionFSM.scala 20:27]
  assign initialOp_io_text = textReg; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 42:25]
  assign initialOp_io_key = keyReg; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 43:24]
  assign finalOp_io_in_state_0_0 = dataReg_state_0_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_0_1 = dataReg_state_0_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_0_2 = dataReg_state_0_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_0_3 = dataReg_state_0_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_1_0 = dataReg_state_1_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_1_1 = dataReg_state_1_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_1_2 = dataReg_state_1_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_1_3 = dataReg_state_1_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_2_0 = dataReg_state_2_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_2_1 = dataReg_state_2_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_2_2 = dataReg_state_2_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_2_3 = dataReg_state_2_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_3_0 = dataReg_state_3_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_3_1 = dataReg_state_3_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_3_2 = dataReg_state_3_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_state_3_3 = dataReg_state_3_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_0_0 = dataReg_key_0_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_0_1 = dataReg_key_0_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_0_2 = dataReg_key_0_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_0_3 = dataReg_key_0_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_1_0 = dataReg_key_1_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_1_1 = dataReg_key_1_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_1_2 = dataReg_key_1_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_1_3 = dataReg_key_1_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_2_0 = dataReg_key_2_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_2_1 = dataReg_key_2_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_2_2 = dataReg_key_2_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_2_3 = dataReg_key_2_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_3_0 = dataReg_key_3_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_3_1 = dataReg_key_3_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_3_2 = dataReg_key_3_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign finalOp_io_in_key_3_3 = dataReg_key_3_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 58:21]
  assign pe_io_in_state_0_0 = dataReg_state_0_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_0_1 = dataReg_state_0_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_0_2 = dataReg_state_0_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_0_3 = dataReg_state_0_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_1_0 = dataReg_state_1_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_1_1 = dataReg_state_1_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_1_2 = dataReg_state_1_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_1_3 = dataReg_state_1_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_2_0 = dataReg_state_2_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_2_1 = dataReg_state_2_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_2_2 = dataReg_state_2_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_2_3 = dataReg_state_2_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_3_0 = dataReg_state_3_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_3_1 = dataReg_state_3_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_3_2 = dataReg_state_3_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_state_3_3 = dataReg_state_3_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_0_0 = dataReg_key_0_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_0_1 = dataReg_key_0_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_0_2 = dataReg_key_0_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_0_3 = dataReg_key_0_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_1_0 = dataReg_key_1_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_1_1 = dataReg_key_1_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_1_2 = dataReg_key_1_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_1_3 = dataReg_key_1_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_2_0 = dataReg_key_2_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_2_1 = dataReg_key_2_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_2_2 = dataReg_key_2_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_2_3 = dataReg_key_2_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_3_0 = dataReg_key_3_0; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_3_1 = dataReg_key_3_1; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_3_2 = dataReg_key_3_2; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_in_key_3_3 = dataReg_key_3_3; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 49:16]
  assign pe_io_round = roundReg; // @[Conditional.scala 39:67 AES_EncryptionFSM.scala 50:19]
  always @(posedge clock) begin
    if (reset) begin // @[AES_EncryptionFSM.scala 13:25]
      stateReg <= 3'h0; // @[AES_EncryptionFSM.scala 13:25]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io_in_valid) begin // @[AES_EncryptionFSM.scala 35:25]
        stateReg <= 3'h1; // @[AES_EncryptionFSM.scala 38:18]
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      stateReg <= 3'h2; // @[AES_EncryptionFSM.scala 46:16]
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      stateReg <= _GEN_3;
    end else begin
      stateReg <= _GEN_40;
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 14:25]
      roundReg <= 4'h0; // @[AES_EncryptionFSM.scala 14:25]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        roundReg <= 4'h0; // @[AES_EncryptionFSM.scala 45:16]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        roundReg <= _T_6; // @[AES_EncryptionFSM.scala 52:16]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 15:24]
      textReg <= 128'h0; // @[AES_EncryptionFSM.scala 15:24]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io_in_valid) begin // @[AES_EncryptionFSM.scala 35:25]
        textReg <= io_in_bits_text; // @[AES_EncryptionFSM.scala 36:17]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 16:23]
      keyReg <= 128'h0; // @[AES_EncryptionFSM.scala 16:23]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io_in_valid) begin // @[AES_EncryptionFSM.scala 35:25]
        keyReg <= io_in_bits_key; // @[AES_EncryptionFSM.scala 37:16]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_0_0 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_0_0 <= initialOp_io_out_state_0_0; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_0_0 <= pe_io_out_state_0_0; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_0_1 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_0_1 <= initialOp_io_out_state_0_1; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_0_1 <= pe_io_out_state_0_1; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_0_2 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_0_2 <= initialOp_io_out_state_0_2; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_0_2 <= pe_io_out_state_0_2; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_0_3 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_0_3 <= initialOp_io_out_state_0_3; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_0_3 <= pe_io_out_state_0_3; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_1_0 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_1_0 <= initialOp_io_out_state_1_0; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_1_0 <= pe_io_out_state_1_0; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_1_1 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_1_1 <= initialOp_io_out_state_1_1; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_1_1 <= pe_io_out_state_1_1; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_1_2 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_1_2 <= initialOp_io_out_state_1_2; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_1_2 <= pe_io_out_state_1_2; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_1_3 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_1_3 <= initialOp_io_out_state_1_3; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_1_3 <= pe_io_out_state_1_3; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_2_0 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_2_0 <= initialOp_io_out_state_2_0; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_2_0 <= pe_io_out_state_2_0; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_2_1 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_2_1 <= initialOp_io_out_state_2_1; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_2_1 <= pe_io_out_state_2_1; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_2_2 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_2_2 <= initialOp_io_out_state_2_2; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_2_2 <= pe_io_out_state_2_2; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_2_3 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_2_3 <= initialOp_io_out_state_2_3; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_2_3 <= pe_io_out_state_2_3; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_3_0 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_3_0 <= initialOp_io_out_state_3_0; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_3_0 <= pe_io_out_state_3_0; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_3_1 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_3_1 <= initialOp_io_out_state_3_1; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_3_1 <= pe_io_out_state_3_1; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_3_2 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_3_2 <= initialOp_io_out_state_3_2; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_3_2 <= pe_io_out_state_3_2; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_state_3_3 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_state_3_3 <= initialOp_io_out_state_3_3; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_state_3_3 <= pe_io_out_state_3_3; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_0_0 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_0_0 <= initialOp_io_out_key_0_0; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_0_0 <= pe_io_out_key_0_0; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_0_1 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_0_1 <= initialOp_io_out_key_0_1; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_0_1 <= pe_io_out_key_0_1; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_0_2 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_0_2 <= initialOp_io_out_key_0_2; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_0_2 <= pe_io_out_key_0_2; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_0_3 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_0_3 <= initialOp_io_out_key_0_3; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_0_3 <= pe_io_out_key_0_3; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_1_0 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_1_0 <= initialOp_io_out_key_1_0; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_1_0 <= pe_io_out_key_1_0; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_1_1 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_1_1 <= initialOp_io_out_key_1_1; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_1_1 <= pe_io_out_key_1_1; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_1_2 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_1_2 <= initialOp_io_out_key_1_2; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_1_2 <= pe_io_out_key_1_2; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_1_3 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_1_3 <= initialOp_io_out_key_1_3; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_1_3 <= pe_io_out_key_1_3; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_2_0 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_2_0 <= initialOp_io_out_key_2_0; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_2_0 <= pe_io_out_key_2_0; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_2_1 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_2_1 <= initialOp_io_out_key_2_1; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_2_1 <= pe_io_out_key_2_1; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_2_2 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_2_2 <= initialOp_io_out_key_2_2; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_2_2 <= pe_io_out_key_2_2; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_2_3 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_2_3 <= initialOp_io_out_key_2_3; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_2_3 <= pe_io_out_key_2_3; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_3_0 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_3_0 <= initialOp_io_out_key_3_0; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_3_0 <= pe_io_out_key_3_0; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_3_1 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_3_1 <= initialOp_io_out_key_3_1; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_3_1 <= pe_io_out_key_3_1; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_3_2 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_3_2 <= initialOp_io_out_key_3_2; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_3_2 <= pe_io_out_key_3_2; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 17:24]
      dataReg_key_3_3 <= 8'h0; // @[AES_EncryptionFSM.scala 17:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_key_3_3 <= initialOp_io_out_key_3_3; // @[AES_EncryptionFSM.scala 44:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_key_3_3 <= pe_io_out_key_3_3; // @[AES_EncryptionFSM.scala 51:15]
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 18:27]
      resultsReg_text <= 128'h0; // @[AES_EncryptionFSM.scala 18:27]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (!(_T_3)) begin // @[Conditional.scala 39:67]
        if (!(_T_4)) begin // @[Conditional.scala 39:67]
          resultsReg_text <= _GEN_39;
        end
      end
    end
    if (reset) begin // @[AES_EncryptionFSM.scala 18:27]
      resultsReg_key <= 128'h0; // @[AES_EncryptionFSM.scala 18:27]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (!(_T_3)) begin // @[Conditional.scala 39:67]
        if (!(_T_4)) begin // @[Conditional.scala 39:67]
          resultsReg_key <= _GEN_38;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  roundReg = _RAND_1[3:0];
  _RAND_2 = {4{`RANDOM}};
  textReg = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  keyReg = _RAND_3[127:0];
  _RAND_4 = {1{`RANDOM}};
  dataReg_state_0_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  dataReg_state_0_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  dataReg_state_0_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  dataReg_state_0_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  dataReg_state_1_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  dataReg_state_1_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  dataReg_state_1_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  dataReg_state_1_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  dataReg_state_2_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  dataReg_state_2_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  dataReg_state_2_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  dataReg_state_2_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  dataReg_state_3_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  dataReg_state_3_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  dataReg_state_3_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  dataReg_state_3_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  dataReg_key_0_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  dataReg_key_0_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  dataReg_key_0_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  dataReg_key_0_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  dataReg_key_1_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  dataReg_key_1_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  dataReg_key_1_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  dataReg_key_1_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  dataReg_key_2_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  dataReg_key_2_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  dataReg_key_2_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  dataReg_key_2_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  dataReg_key_3_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  dataReg_key_3_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  dataReg_key_3_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  dataReg_key_3_3 = _RAND_35[7:0];
  _RAND_36 = {4{`RANDOM}};
  resultsReg_text = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  resultsReg_key = _RAND_37[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
