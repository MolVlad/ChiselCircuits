module AES_InitialOperation(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits_text,
  input  [127:0] io_in_bits_key,
  input          io_out_ready,
  output         io_out_valid,
  output [7:0]   io_out_bits_state_0_0,
  output [7:0]   io_out_bits_state_0_1,
  output [7:0]   io_out_bits_state_0_2,
  output [7:0]   io_out_bits_state_0_3,
  output [7:0]   io_out_bits_state_1_0,
  output [7:0]   io_out_bits_state_1_1,
  output [7:0]   io_out_bits_state_1_2,
  output [7:0]   io_out_bits_state_1_3,
  output [7:0]   io_out_bits_state_2_0,
  output [7:0]   io_out_bits_state_2_1,
  output [7:0]   io_out_bits_state_2_2,
  output [7:0]   io_out_bits_state_2_3,
  output [7:0]   io_out_bits_state_3_0,
  output [7:0]   io_out_bits_state_3_1,
  output [7:0]   io_out_bits_state_3_2,
  output [7:0]   io_out_bits_state_3_3,
  output [7:0]   io_out_bits_key_0_0,
  output [7:0]   io_out_bits_key_0_1,
  output [7:0]   io_out_bits_key_0_2,
  output [7:0]   io_out_bits_key_0_3,
  output [7:0]   io_out_bits_key_1_0,
  output [7:0]   io_out_bits_key_1_1,
  output [7:0]   io_out_bits_key_1_2,
  output [7:0]   io_out_bits_key_1_3,
  output [7:0]   io_out_bits_key_2_0,
  output [7:0]   io_out_bits_key_2_1,
  output [7:0]   io_out_bits_key_2_2,
  output [7:0]   io_out_bits_key_2_3,
  output [7:0]   io_out_bits_key_3_0,
  output [7:0]   io_out_bits_key_3_1,
  output [7:0]   io_out_bits_key_3_2,
  output [7:0]   io_out_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] data_0_text; // @[AES_PipelinedElasticBuffer.scala 58:21]
  reg [127:0] data_0_key; // @[AES_PipelinedElasticBuffer.scala 58:21]
  reg [127:0] data_1_text; // @[AES_PipelinedElasticBuffer.scala 58:21]
  reg [127:0] data_1_key; // @[AES_PipelinedElasticBuffer.scala 58:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 59:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 60:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 61:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 61:21]
  wire [127:0] input_text = head ? data_1_text : data_0_text; // @[AES_PipelinedElasticBuffer.scala 66:9 AES_PipelinedElasticBuffer.scala 66:9]
  wire [127:0] input_key = head ? data_1_key : data_0_key; // @[AES_PipelinedElasticBuffer.scala 66:9 AES_PipelinedElasticBuffer.scala 66:9]
  wire  _GEN_5 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 69:23 AES_PipelinedElasticBuffer.scala 69:23]
  wire  _GEN_26 = ~tail; // @[AES_PipelinedElasticBuffer.scala 70:16 AES_PipelinedElasticBuffer.scala 70:16 AES_PipelinedElasticBuffer.scala 61:21]
  wire  _GEN_6 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 70:16 AES_PipelinedElasticBuffer.scala 70:16 AES_PipelinedElasticBuffer.scala 61:21]
  wire  _GEN_7 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 70:16 AES_PipelinedElasticBuffer.scala 70:16 AES_PipelinedElasticBuffer.scala 61:21]
  wire  _GEN_12 = io_in_valid & ~_GEN_5 ? _GEN_6 : full_0; // @[AES_PipelinedElasticBuffer.scala 69:36 AES_PipelinedElasticBuffer.scala 61:21]
  wire  _GEN_13 = io_in_valid & ~_GEN_5 ? _GEN_7 : full_1; // @[AES_PipelinedElasticBuffer.scala 69:36 AES_PipelinedElasticBuffer.scala 61:21]
  wire  _GEN_20 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 76:21 AES_PipelinedElasticBuffer.scala 76:21]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 63:18]
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 64:27]
  assign io_out_bits_state_0_0 = input_text[127:120]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_0_1 = input_text[119:112]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_0_2 = input_text[111:104]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_0_3 = input_text[103:96]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_1_0 = input_text[95:88]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_1_1 = input_text[87:80]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_1_2 = input_text[79:72]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_1_3 = input_text[71:64]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_2_0 = input_text[63:56]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_2_1 = input_text[55:48]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_2_2 = input_text[47:40]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_2_3 = input_text[39:32]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_3_0 = input_text[31:24]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_3_1 = input_text[23:16]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_3_2 = input_text[15:8]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_state_3_3 = input_text[7:0]; // @[AES_PipelinedElasticBuffer.scala 84:43]
  assign io_out_bits_key_0_0 = input_key[127:120]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_0_1 = input_key[119:112]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_0_2 = input_key[111:104]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_0_3 = input_key[103:96]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_1_0 = input_key[95:88]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_1_1 = input_key[87:80]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_1_2 = input_key[79:72]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_1_3 = input_key[71:64]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_2_0 = input_key[63:56]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_2_1 = input_key[55:48]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_2_2 = input_key[47:40]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_2_3 = input_key[39:32]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_3_0 = input_key[31:24]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_3_1 = input_key[23:16]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_3_2 = input_key[15:8]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  assign io_out_bits_key_3_3 = input_key[7:0]; // @[AES_PipelinedElasticBuffer.scala 85:40]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 58:21]
      data_0_text <= 128'h0; // @[AES_PipelinedElasticBuffer.scala 58:21]
    end else if (io_in_valid & ~_GEN_5) begin // @[AES_PipelinedElasticBuffer.scala 69:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 71:16]
        data_0_text <= io_in_bits_text; // @[AES_PipelinedElasticBuffer.scala 71:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 58:21]
      data_0_key <= 128'h0; // @[AES_PipelinedElasticBuffer.scala 58:21]
    end else if (io_in_valid & ~_GEN_5) begin // @[AES_PipelinedElasticBuffer.scala 69:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 71:16]
        data_0_key <= io_in_bits_key; // @[AES_PipelinedElasticBuffer.scala 71:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 58:21]
      data_1_text <= 128'h0; // @[AES_PipelinedElasticBuffer.scala 58:21]
    end else if (io_in_valid & ~_GEN_5) begin // @[AES_PipelinedElasticBuffer.scala 69:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 71:16]
        data_1_text <= io_in_bits_text; // @[AES_PipelinedElasticBuffer.scala 71:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 58:21]
      data_1_key <= 128'h0; // @[AES_PipelinedElasticBuffer.scala 58:21]
    end else if (io_in_valid & ~_GEN_5) begin // @[AES_PipelinedElasticBuffer.scala 69:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 71:16]
        data_1_key <= io_in_bits_key; // @[AES_PipelinedElasticBuffer.scala 71:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 59:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 59:21]
    end else if (io_out_ready & _GEN_20) begin // @[AES_PipelinedElasticBuffer.scala 76:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 78:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 60:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 60:21]
    end else if (io_in_valid & ~_GEN_5) begin // @[AES_PipelinedElasticBuffer.scala 69:36]
      tail <= _GEN_26; // @[AES_PipelinedElasticBuffer.scala 72:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 61:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 61:21]
    end else if (io_out_ready & _GEN_20) begin // @[AES_PipelinedElasticBuffer.scala 76:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 77:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 77:16]
      end else begin
        full_0 <= _GEN_12;
      end
    end else begin
      full_0 <= _GEN_12;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 61:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 61:21]
    end else if (io_out_ready & _GEN_20) begin // @[AES_PipelinedElasticBuffer.scala 76:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 77:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 77:16]
      end else begin
        full_1 <= _GEN_13;
      end
    end else begin
      full_1 <= _GEN_13;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  data_0_text = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  data_0_key = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  data_1_text = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  data_1_key = _RAND_3[127:0];
  _RAND_4 = {1{`RANDOM}};
  head = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tail = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  full_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  full_1 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_FinalOperation(
  input          clock,
  input          reset,
  input          io_out_ready,
  output         io_out_valid,
  output [127:0] io_out_bits_text,
  output [127:0] io_out_bits_key,
  output         io_in_ready,
  input          io_in_valid,
  input  [7:0]   io_in_bits_state_0_0,
  input  [7:0]   io_in_bits_state_0_1,
  input  [7:0]   io_in_bits_state_0_2,
  input  [7:0]   io_in_bits_state_0_3,
  input  [7:0]   io_in_bits_state_1_0,
  input  [7:0]   io_in_bits_state_1_1,
  input  [7:0]   io_in_bits_state_1_2,
  input  [7:0]   io_in_bits_state_1_3,
  input  [7:0]   io_in_bits_state_2_0,
  input  [7:0]   io_in_bits_state_2_1,
  input  [7:0]   io_in_bits_state_2_2,
  input  [7:0]   io_in_bits_state_2_3,
  input  [7:0]   io_in_bits_state_3_0,
  input  [7:0]   io_in_bits_state_3_1,
  input  [7:0]   io_in_bits_state_3_2,
  input  [7:0]   io_in_bits_state_3_3,
  input  [7:0]   io_in_bits_key_0_0,
  input  [7:0]   io_in_bits_key_0_1,
  input  [7:0]   io_in_bits_key_0_2,
  input  [7:0]   io_in_bits_key_0_3,
  input  [7:0]   io_in_bits_key_1_0,
  input  [7:0]   io_in_bits_key_1_1,
  input  [7:0]   io_in_bits_key_1_2,
  input  [7:0]   io_in_bits_key_1_3,
  input  [7:0]   io_in_bits_key_2_0,
  input  [7:0]   io_in_bits_key_2_1,
  input  [7:0]   io_in_bits_key_2_2,
  input  [7:0]   io_in_bits_key_2_3,
  input  [7:0]   io_in_bits_key_3_0,
  input  [7:0]   io_in_bits_key_3_1,
  input  [7:0]   io_in_bits_key_3_2,
  input  [7:0]   io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 98:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 99:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 100:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 101:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 101:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 106:9 AES_PipelinedElasticBuffer.scala 106:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 109:23 AES_PipelinedElasticBuffer.scala 109:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 110:16 AES_PipelinedElasticBuffer.scala 110:16 AES_PipelinedElasticBuffer.scala 101:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 110:16 AES_PipelinedElasticBuffer.scala 110:16 AES_PipelinedElasticBuffer.scala 101:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 110:16 AES_PipelinedElasticBuffer.scala 110:16 AES_PipelinedElasticBuffer.scala 101:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 109:36 AES_PipelinedElasticBuffer.scala 101:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 109:36 AES_PipelinedElasticBuffer.scala 101:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 116:21 AES_PipelinedElasticBuffer.scala 116:21]
  wire [7:0] hi_hi_hi_hi = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 122:39]
  wire [7:0] hi_hi_hi_lo = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 122:73]
  wire [7:0] hi_hi_lo_hi = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 123:22]
  wire [7:0] hi_hi_lo_lo = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 123:56]
  wire [7:0] hi_lo_hi_hi = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 124:22]
  wire [7:0] hi_lo_hi_lo = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 124:56]
  wire [7:0] hi_lo_lo_hi = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 125:22]
  wire [7:0] hi_lo_lo_lo = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 125:56]
  wire [7:0] lo_hi_hi_hi = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 126:22]
  wire [7:0] lo_hi_hi_lo = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 126:56]
  wire [7:0] lo_hi_lo_hi = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 127:22]
  wire [7:0] lo_hi_lo_lo = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 127:56]
  wire [7:0] lo_lo_hi_hi = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 128:22]
  wire [7:0] lo_lo_hi_lo = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 128:56]
  wire [7:0] lo_lo_lo_hi = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 129:22]
  wire [7:0] lo_lo_lo_lo = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 129:56]
  wire [63:0] lo = {lo_hi_hi_hi,lo_hi_hi_lo,lo_hi_lo_hi,lo_hi_lo_lo,lo_lo_hi_hi,lo_lo_hi_lo,lo_lo_lo_hi,lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] hi = {hi_hi_hi_hi,hi_hi_hi_lo,hi_hi_lo_hi,hi_hi_lo_lo,hi_lo_hi_hi,hi_lo_hi_lo,hi_lo_lo_hi,hi_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] lo_1 = {input_key_2_0,input_key_2_1,input_key_2_2,input_key_2_3,input_key_3_0,input_key_3_1,input_key_3_2,
    input_key_3_3}; // @[Cat.scala 30:58]
  wire [63:0] hi_1 = {input_key_0_0,input_key_0_1,input_key_0_2,input_key_0_3,input_key_1_0,input_key_1_1,input_key_1_2,
    input_key_1_3}; // @[Cat.scala 30:58]
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 104:27]
  assign io_out_bits_text = {hi,lo}; // @[Cat.scala 30:58]
  assign io_out_bits_key = {hi_1,lo_1}; // @[Cat.scala 30:58]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 103:18]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 98:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 98:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 111:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 111:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 99:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 99:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 118:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 100:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 100:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 109:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 112:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 101:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 101:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 117:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 117:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 101:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 101:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 117:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 117:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_XOR(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  assign io_out_state_0_0 = io_in_state_0_0 ^ io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_0_1 = io_in_state_0_1 ^ io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_0_2 = io_in_state_0_2 ^ io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_0_3 = io_in_state_0_3 ^ io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_1_0 = io_in_state_1_0 ^ io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_1_1 = io_in_state_1_1 ^ io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_1_2 = io_in_state_1_2 ^ io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_1_3 = io_in_state_1_3 ^ io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_2_0 = io_in_state_2_0 ^ io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_2_1 = io_in_state_2_1 ^ io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_2_2 = io_in_state_2_2 ^ io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_2_3 = io_in_state_2_3 ^ io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_3_0 = io_in_state_3_0 ^ io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_3_1 = io_in_state_3_1 ^ io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_3_2 = io_in_state_3_2 ^ io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 330:47]
  assign io_out_state_3_3 = io_in_state_3_3 ^ io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 330:47]
endmodule
module AES_S(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _GEN_1 = 4'h0 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h7c : 8'h63; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_2 = 4'h0 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h77 : _GEN_1; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_3 = 4'h0 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h7b : _GEN_2; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_4 = 4'h0 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hf2 : _GEN_3; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_5 = 4'h0 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h6b : _GEN_4; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_6 = 4'h0 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h6f : _GEN_5; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_7 = 4'h0 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hc5 : _GEN_6; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_8 = 4'h0 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h30 : _GEN_7; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_9 = 4'h0 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h1 : _GEN_8; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_10 = 4'h0 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h67 : _GEN_9; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_11 = 4'h0 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h2b : _GEN_10; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_12 = 4'h0 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hfe : _GEN_11; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_13 = 4'h0 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hd7 : _GEN_12; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_14 = 4'h0 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hab : _GEN_13; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_15 = 4'h0 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h76 : _GEN_14; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_16 = 4'h1 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hca : _GEN_15; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_17 = 4'h1 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h82 : _GEN_16; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_18 = 4'h1 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'hc9 : _GEN_17; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_19 = 4'h1 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h7d : _GEN_18; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_20 = 4'h1 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hfa : _GEN_19; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_21 = 4'h1 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h59 : _GEN_20; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_22 = 4'h1 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h47 : _GEN_21; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_23 = 4'h1 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hf0 : _GEN_22; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_24 = 4'h1 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'had : _GEN_23; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_25 = 4'h1 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hd4 : _GEN_24; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_26 = 4'h1 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'ha2 : _GEN_25; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_27 = 4'h1 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'haf : _GEN_26; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_28 = 4'h1 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h9c : _GEN_27; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_29 = 4'h1 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'ha4 : _GEN_28; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_30 = 4'h1 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h72 : _GEN_29; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_31 = 4'h1 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hc0 : _GEN_30; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_32 = 4'h2 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hb7 : _GEN_31; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_33 = 4'h2 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hfd : _GEN_32; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_34 = 4'h2 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h93 : _GEN_33; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_35 = 4'h2 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h26 : _GEN_34; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_36 = 4'h2 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h36 : _GEN_35; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_37 = 4'h2 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h3f : _GEN_36; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_38 = 4'h2 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hf7 : _GEN_37; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_39 = 4'h2 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hcc : _GEN_38; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_40 = 4'h2 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h34 : _GEN_39; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_41 = 4'h2 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'ha5 : _GEN_40; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_42 = 4'h2 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'he5 : _GEN_41; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_43 = 4'h2 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hf1 : _GEN_42; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_44 = 4'h2 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h71 : _GEN_43; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_45 = 4'h2 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hd8 : _GEN_44; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_46 = 4'h2 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h31 : _GEN_45; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_47 = 4'h2 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h15 : _GEN_46; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_48 = 4'h3 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h4 : _GEN_47; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_49 = 4'h3 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hc7 : _GEN_48; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_50 = 4'h3 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h23 : _GEN_49; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_51 = 4'h3 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hc3 : _GEN_50; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_52 = 4'h3 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h18 : _GEN_51; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_53 = 4'h3 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h96 : _GEN_52; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_54 = 4'h3 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h5 : _GEN_53; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_55 = 4'h3 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h9a : _GEN_54; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_56 = 4'h3 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h7 : _GEN_55; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_57 = 4'h3 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h12 : _GEN_56; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_58 = 4'h3 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h80 : _GEN_57; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_59 = 4'h3 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'he2 : _GEN_58; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_60 = 4'h3 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'heb : _GEN_59; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_61 = 4'h3 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h27 : _GEN_60; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_62 = 4'h3 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hb2 : _GEN_61; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_63 = 4'h3 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h75 : _GEN_62; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_64 = 4'h4 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h9 : _GEN_63; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_65 = 4'h4 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h83 : _GEN_64; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_66 = 4'h4 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h2c : _GEN_65; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_67 = 4'h4 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h1a : _GEN_66; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_68 = 4'h4 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h1b : _GEN_67; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_69 = 4'h4 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h6e : _GEN_68; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_70 = 4'h4 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h5a : _GEN_69; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_71 = 4'h4 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'ha0 : _GEN_70; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_72 = 4'h4 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h52 : _GEN_71; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_73 = 4'h4 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h3b : _GEN_72; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_74 = 4'h4 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hd6 : _GEN_73; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_75 = 4'h4 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hb3 : _GEN_74; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_76 = 4'h4 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h29 : _GEN_75; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_77 = 4'h4 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'he3 : _GEN_76; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_78 = 4'h4 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h2f : _GEN_77; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_79 = 4'h4 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h84 : _GEN_78; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_80 = 4'h5 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h53 : _GEN_79; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_81 = 4'h5 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hd1 : _GEN_80; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_82 = 4'h5 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h0 : _GEN_81; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_83 = 4'h5 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hed : _GEN_82; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_84 = 4'h5 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h20 : _GEN_83; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_85 = 4'h5 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hfc : _GEN_84; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_86 = 4'h5 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hb1 : _GEN_85; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_87 = 4'h5 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h5b : _GEN_86; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_88 = 4'h5 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h6a : _GEN_87; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_89 = 4'h5 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hcb : _GEN_88; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_90 = 4'h5 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hbe : _GEN_89; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_91 = 4'h5 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h39 : _GEN_90; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_92 = 4'h5 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h4a : _GEN_91; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_93 = 4'h5 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h4c : _GEN_92; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_94 = 4'h5 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h58 : _GEN_93; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_95 = 4'h5 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hcf : _GEN_94; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_96 = 4'h6 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hd0 : _GEN_95; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_97 = 4'h6 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hef : _GEN_96; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_98 = 4'h6 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'haa : _GEN_97; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_99 = 4'h6 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hfb : _GEN_98; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_100 = 4'h6 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h43 : _GEN_99; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_101 = 4'h6 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h4d : _GEN_100; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_102 = 4'h6 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h33 : _GEN_101; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_103 = 4'h6 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h85 : _GEN_102; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_104 = 4'h6 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h45 : _GEN_103; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_105 = 4'h6 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hf9 : _GEN_104; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_106 = 4'h6 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h2 : _GEN_105; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_107 = 4'h6 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h7f : _GEN_106; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_108 = 4'h6 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h50 : _GEN_107; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_109 = 4'h6 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h3c : _GEN_108; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_110 = 4'h6 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h9f : _GEN_109; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_111 = 4'h6 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'ha8 : _GEN_110; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_112 = 4'h7 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h51 : _GEN_111; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_113 = 4'h7 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'ha3 : _GEN_112; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_114 = 4'h7 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h40 : _GEN_113; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_115 = 4'h7 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h8f : _GEN_114; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_116 = 4'h7 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h92 : _GEN_115; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_117 = 4'h7 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h9d : _GEN_116; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_118 = 4'h7 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h38 : _GEN_117; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_119 = 4'h7 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hf5 : _GEN_118; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_120 = 4'h7 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hbc : _GEN_119; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_121 = 4'h7 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hb6 : _GEN_120; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_122 = 4'h7 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hda : _GEN_121; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_123 = 4'h7 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h21 : _GEN_122; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_124 = 4'h7 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h10 : _GEN_123; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_125 = 4'h7 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hff : _GEN_124; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_126 = 4'h7 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hf3 : _GEN_125; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_127 = 4'h7 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hd2 : _GEN_126; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_128 = 4'h8 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hcd : _GEN_127; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_129 = 4'h8 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hc : _GEN_128; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_130 = 4'h8 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h13 : _GEN_129; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_131 = 4'h8 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hec : _GEN_130; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_132 = 4'h8 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h5f : _GEN_131; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_133 = 4'h8 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h97 : _GEN_132; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_134 = 4'h8 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h44 : _GEN_133; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_135 = 4'h8 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h17 : _GEN_134; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_136 = 4'h8 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hc4 : _GEN_135; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_137 = 4'h8 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'ha7 : _GEN_136; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_138 = 4'h8 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h7e : _GEN_137; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_139 = 4'h8 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h3d : _GEN_138; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_140 = 4'h8 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h64 : _GEN_139; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_141 = 4'h8 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h5d : _GEN_140; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_142 = 4'h8 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h19 : _GEN_141; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_143 = 4'h8 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h73 : _GEN_142; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_144 = 4'h9 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h60 : _GEN_143; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_145 = 4'h9 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h81 : _GEN_144; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_146 = 4'h9 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h4f : _GEN_145; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_147 = 4'h9 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hdc : _GEN_146; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_148 = 4'h9 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h22 : _GEN_147; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_149 = 4'h9 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h2a : _GEN_148; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_150 = 4'h9 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h90 : _GEN_149; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_151 = 4'h9 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h88 : _GEN_150; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_152 = 4'h9 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h46 : _GEN_151; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_153 = 4'h9 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hee : _GEN_152; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_154 = 4'h9 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hb8 : _GEN_153; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_155 = 4'h9 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h14 : _GEN_154; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_156 = 4'h9 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hde : _GEN_155; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_157 = 4'h9 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h5e : _GEN_156; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_158 = 4'h9 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hb : _GEN_157; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_159 = 4'h9 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hdb : _GEN_158; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_160 = 4'ha == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'he0 : _GEN_159; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_161 = 4'ha == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h32 : _GEN_160; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_162 = 4'ha == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h3a : _GEN_161; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_163 = 4'ha == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'ha : _GEN_162; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_164 = 4'ha == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h49 : _GEN_163; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_165 = 4'ha == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h6 : _GEN_164; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_166 = 4'ha == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h24 : _GEN_165; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_167 = 4'ha == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h5c : _GEN_166; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_168 = 4'ha == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hc2 : _GEN_167; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_169 = 4'ha == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hd3 : _GEN_168; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_170 = 4'ha == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hac : _GEN_169; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_171 = 4'ha == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h62 : _GEN_170; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_172 = 4'ha == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h91 : _GEN_171; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_173 = 4'ha == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h95 : _GEN_172; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_174 = 4'ha == io_in[7:4] & 4'he == io_in[3:0] ? 8'he4 : _GEN_173; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_175 = 4'ha == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h79 : _GEN_174; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_176 = 4'hb == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'he7 : _GEN_175; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_177 = 4'hb == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hc8 : _GEN_176; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_178 = 4'hb == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h37 : _GEN_177; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_179 = 4'hb == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h6d : _GEN_178; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_180 = 4'hb == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h8d : _GEN_179; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_181 = 4'hb == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hd5 : _GEN_180; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_182 = 4'hb == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h4e : _GEN_181; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_183 = 4'hb == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'ha9 : _GEN_182; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_184 = 4'hb == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h6c : _GEN_183; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_185 = 4'hb == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h56 : _GEN_184; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_186 = 4'hb == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hf4 : _GEN_185; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_187 = 4'hb == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hea : _GEN_186; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_188 = 4'hb == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h65 : _GEN_187; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_189 = 4'hb == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h7a : _GEN_188; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_190 = 4'hb == io_in[7:4] & 4'he == io_in[3:0] ? 8'hae : _GEN_189; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_191 = 4'hb == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h8 : _GEN_190; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_192 = 4'hc == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hba : _GEN_191; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_193 = 4'hc == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h78 : _GEN_192; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_194 = 4'hc == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h25 : _GEN_193; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_195 = 4'hc == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h2e : _GEN_194; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_196 = 4'hc == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h1c : _GEN_195; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_197 = 4'hc == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'ha6 : _GEN_196; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_198 = 4'hc == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hb4 : _GEN_197; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_199 = 4'hc == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hc6 : _GEN_198; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_200 = 4'hc == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'he8 : _GEN_199; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_201 = 4'hc == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hdd : _GEN_200; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_202 = 4'hc == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h74 : _GEN_201; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_203 = 4'hc == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h1f : _GEN_202; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_204 = 4'hc == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h4b : _GEN_203; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_205 = 4'hc == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hbd : _GEN_204; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_206 = 4'hc == io_in[7:4] & 4'he == io_in[3:0] ? 8'h8b : _GEN_205; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_207 = 4'hc == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h8a : _GEN_206; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_208 = 4'hd == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h70 : _GEN_207; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_209 = 4'hd == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h3e : _GEN_208; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_210 = 4'hd == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'hb5 : _GEN_209; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_211 = 4'hd == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h66 : _GEN_210; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_212 = 4'hd == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h48 : _GEN_211; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_213 = 4'hd == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h3 : _GEN_212; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_214 = 4'hd == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hf6 : _GEN_213; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_215 = 4'hd == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'he : _GEN_214; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_216 = 4'hd == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h61 : _GEN_215; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_217 = 4'hd == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h35 : _GEN_216; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_218 = 4'hd == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h57 : _GEN_217; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_219 = 4'hd == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hb9 : _GEN_218; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_220 = 4'hd == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h86 : _GEN_219; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_221 = 4'hd == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hc1 : _GEN_220; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_222 = 4'hd == io_in[7:4] & 4'he == io_in[3:0] ? 8'h1d : _GEN_221; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_223 = 4'hd == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h9e : _GEN_222; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_224 = 4'he == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'he1 : _GEN_223; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_225 = 4'he == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hf8 : _GEN_224; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_226 = 4'he == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h98 : _GEN_225; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_227 = 4'he == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h11 : _GEN_226; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_228 = 4'he == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h69 : _GEN_227; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_229 = 4'he == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hd9 : _GEN_228; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_230 = 4'he == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h8e : _GEN_229; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_231 = 4'he == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h94 : _GEN_230; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_232 = 4'he == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h9b : _GEN_231; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_233 = 4'he == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h1e : _GEN_232; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_234 = 4'he == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h87 : _GEN_233; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_235 = 4'he == io_in[7:4] & 4'hb == io_in[3:0] ? 8'he9 : _GEN_234; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_236 = 4'he == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hce : _GEN_235; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_237 = 4'he == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h55 : _GEN_236; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_238 = 4'he == io_in[7:4] & 4'he == io_in[3:0] ? 8'h28 : _GEN_237; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_239 = 4'he == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hdf : _GEN_238; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_240 = 4'hf == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h8c : _GEN_239; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_241 = 4'hf == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'ha1 : _GEN_240; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_242 = 4'hf == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h89 : _GEN_241; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_243 = 4'hf == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hd : _GEN_242; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_244 = 4'hf == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hbf : _GEN_243; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_245 = 4'hf == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'he6 : _GEN_244; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_246 = 4'hf == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h42 : _GEN_245; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_247 = 4'hf == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h68 : _GEN_246; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_248 = 4'hf == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h41 : _GEN_247; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_249 = 4'hf == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h99 : _GEN_248; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_250 = 4'hf == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h2d : _GEN_249; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_251 = 4'hf == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hf : _GEN_250; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_252 = 4'hf == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hb0 : _GEN_251; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_253 = 4'hf == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h54 : _GEN_252; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  wire [7:0] _GEN_254 = 4'hf == io_in[7:4] & 4'he == io_in[3:0] ? 8'hbb : _GEN_253; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
  assign io_out = 4'hf == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h16 : _GEN_254; // @[AES_PipelinedElasticBuffer.scala 742:10 AES_PipelinedElasticBuffer.scala 742:10]
endmodule
module AES_SubBytes(
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3
);
  wire [7:0] PEs_0_0_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_0_0_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_0_1_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_0_1_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_0_2_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_0_2_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_0_3_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_0_3_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_1_0_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_1_0_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_1_1_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_1_1_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_1_2_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_1_2_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_1_3_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_1_3_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_2_0_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_2_0_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_2_1_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_2_1_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_2_2_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_2_2_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_2_3_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_2_3_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_3_0_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_3_0_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_3_1_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_3_1_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_3_2_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_3_2_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_3_3_io_in; // @[AES_PipelinedElasticBuffer.scala 665:22]
  wire [7:0] PEs_3_3_io_out; // @[AES_PipelinedElasticBuffer.scala 665:22]
  AES_S PEs_0_0 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_0_0_io_in),
    .io_out(PEs_0_0_io_out)
  );
  AES_S PEs_0_1 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_0_1_io_in),
    .io_out(PEs_0_1_io_out)
  );
  AES_S PEs_0_2 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_0_2_io_in),
    .io_out(PEs_0_2_io_out)
  );
  AES_S PEs_0_3 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_0_3_io_in),
    .io_out(PEs_0_3_io_out)
  );
  AES_S PEs_1_0 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_1_0_io_in),
    .io_out(PEs_1_0_io_out)
  );
  AES_S PEs_1_1 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_1_1_io_in),
    .io_out(PEs_1_1_io_out)
  );
  AES_S PEs_1_2 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_1_2_io_in),
    .io_out(PEs_1_2_io_out)
  );
  AES_S PEs_1_3 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_1_3_io_in),
    .io_out(PEs_1_3_io_out)
  );
  AES_S PEs_2_0 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_2_0_io_in),
    .io_out(PEs_2_0_io_out)
  );
  AES_S PEs_2_1 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_2_1_io_in),
    .io_out(PEs_2_1_io_out)
  );
  AES_S PEs_2_2 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_2_2_io_in),
    .io_out(PEs_2_2_io_out)
  );
  AES_S PEs_2_3 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_2_3_io_in),
    .io_out(PEs_2_3_io_out)
  );
  AES_S PEs_3_0 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_3_0_io_in),
    .io_out(PEs_3_0_io_out)
  );
  AES_S PEs_3_1 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_3_1_io_in),
    .io_out(PEs_3_1_io_out)
  );
  AES_S PEs_3_2 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_3_2_io_in),
    .io_out(PEs_3_2_io_out)
  );
  AES_S PEs_3_3 ( // @[AES_PipelinedElasticBuffer.scala 665:22]
    .io_in(PEs_3_3_io_in),
    .io_out(PEs_3_3_io_out)
  );
  assign PEs_0_0_io_in = io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_0_1_io_in = io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_0_2_io_in = io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_0_3_io_in = io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_1_0_io_in = io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_1_1_io_in = io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_1_2_io_in = io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_1_3_io_in = io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_2_0_io_in = io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_2_1_io_in = io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_2_2_io_in = io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_2_3_io_in = io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_3_0_io_in = io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_3_1_io_in = io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_3_2_io_in = io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 673:25]
  assign PEs_3_3_io_in = io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 673:25]
endmodule
module AES_InvMixColumn(
  input  [7:0] io_in_0,
  input  [7:0] io_in_1,
  input  [7:0] io_in_2,
  input  [7:0] io_in_3,
  output [7:0] io_out_0,
  output [7:0] io_out_1,
  output [7:0] io_out_2,
  output [7:0] io_out_3
);
  wire [7:0] _GEN_1 = 8'h1 == io_in_0 ? 8'he : 8'h0; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_2 = 8'h2 == io_in_0 ? 8'h1c : _GEN_1; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_3 = 8'h3 == io_in_0 ? 8'h12 : _GEN_2; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_4 = 8'h4 == io_in_0 ? 8'h38 : _GEN_3; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_5 = 8'h5 == io_in_0 ? 8'h36 : _GEN_4; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_6 = 8'h6 == io_in_0 ? 8'h24 : _GEN_5; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_7 = 8'h7 == io_in_0 ? 8'h2a : _GEN_6; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_8 = 8'h8 == io_in_0 ? 8'h70 : _GEN_7; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_9 = 8'h9 == io_in_0 ? 8'h7e : _GEN_8; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_10 = 8'ha == io_in_0 ? 8'h6c : _GEN_9; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_11 = 8'hb == io_in_0 ? 8'h62 : _GEN_10; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_12 = 8'hc == io_in_0 ? 8'h48 : _GEN_11; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_13 = 8'hd == io_in_0 ? 8'h46 : _GEN_12; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_14 = 8'he == io_in_0 ? 8'h54 : _GEN_13; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_15 = 8'hf == io_in_0 ? 8'h5a : _GEN_14; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_16 = 8'h10 == io_in_0 ? 8'he0 : _GEN_15; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_17 = 8'h11 == io_in_0 ? 8'hee : _GEN_16; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_18 = 8'h12 == io_in_0 ? 8'hfc : _GEN_17; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_19 = 8'h13 == io_in_0 ? 8'hf2 : _GEN_18; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_20 = 8'h14 == io_in_0 ? 8'hd8 : _GEN_19; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_21 = 8'h15 == io_in_0 ? 8'hd6 : _GEN_20; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_22 = 8'h16 == io_in_0 ? 8'hc4 : _GEN_21; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_23 = 8'h17 == io_in_0 ? 8'hca : _GEN_22; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_24 = 8'h18 == io_in_0 ? 8'h90 : _GEN_23; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_25 = 8'h19 == io_in_0 ? 8'h9e : _GEN_24; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_26 = 8'h1a == io_in_0 ? 8'h8c : _GEN_25; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_27 = 8'h1b == io_in_0 ? 8'h82 : _GEN_26; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_28 = 8'h1c == io_in_0 ? 8'ha8 : _GEN_27; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_29 = 8'h1d == io_in_0 ? 8'ha6 : _GEN_28; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_30 = 8'h1e == io_in_0 ? 8'hb4 : _GEN_29; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_31 = 8'h1f == io_in_0 ? 8'hba : _GEN_30; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_32 = 8'h20 == io_in_0 ? 8'hdb : _GEN_31; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_33 = 8'h21 == io_in_0 ? 8'hd5 : _GEN_32; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_34 = 8'h22 == io_in_0 ? 8'hc7 : _GEN_33; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_35 = 8'h23 == io_in_0 ? 8'hc9 : _GEN_34; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_36 = 8'h24 == io_in_0 ? 8'he3 : _GEN_35; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_37 = 8'h25 == io_in_0 ? 8'hed : _GEN_36; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_38 = 8'h26 == io_in_0 ? 8'hff : _GEN_37; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_39 = 8'h27 == io_in_0 ? 8'hf1 : _GEN_38; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_40 = 8'h28 == io_in_0 ? 8'hab : _GEN_39; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_41 = 8'h29 == io_in_0 ? 8'ha5 : _GEN_40; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_42 = 8'h2a == io_in_0 ? 8'hb7 : _GEN_41; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_43 = 8'h2b == io_in_0 ? 8'hb9 : _GEN_42; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_44 = 8'h2c == io_in_0 ? 8'h93 : _GEN_43; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_45 = 8'h2d == io_in_0 ? 8'h9d : _GEN_44; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_46 = 8'h2e == io_in_0 ? 8'h8f : _GEN_45; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_47 = 8'h2f == io_in_0 ? 8'h81 : _GEN_46; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_48 = 8'h30 == io_in_0 ? 8'h3b : _GEN_47; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_49 = 8'h31 == io_in_0 ? 8'h35 : _GEN_48; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_50 = 8'h32 == io_in_0 ? 8'h27 : _GEN_49; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_51 = 8'h33 == io_in_0 ? 8'h29 : _GEN_50; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_52 = 8'h34 == io_in_0 ? 8'h3 : _GEN_51; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_53 = 8'h35 == io_in_0 ? 8'hd : _GEN_52; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_54 = 8'h36 == io_in_0 ? 8'h1f : _GEN_53; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_55 = 8'h37 == io_in_0 ? 8'h11 : _GEN_54; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_56 = 8'h38 == io_in_0 ? 8'h4b : _GEN_55; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_57 = 8'h39 == io_in_0 ? 8'h45 : _GEN_56; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_58 = 8'h3a == io_in_0 ? 8'h57 : _GEN_57; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_59 = 8'h3b == io_in_0 ? 8'h59 : _GEN_58; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_60 = 8'h3c == io_in_0 ? 8'h73 : _GEN_59; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_61 = 8'h3d == io_in_0 ? 8'h7d : _GEN_60; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_62 = 8'h3e == io_in_0 ? 8'h6f : _GEN_61; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_63 = 8'h3f == io_in_0 ? 8'h61 : _GEN_62; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_64 = 8'h40 == io_in_0 ? 8'had : _GEN_63; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_65 = 8'h41 == io_in_0 ? 8'ha3 : _GEN_64; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_66 = 8'h42 == io_in_0 ? 8'hb1 : _GEN_65; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_67 = 8'h43 == io_in_0 ? 8'hbf : _GEN_66; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_68 = 8'h44 == io_in_0 ? 8'h95 : _GEN_67; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_69 = 8'h45 == io_in_0 ? 8'h9b : _GEN_68; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_70 = 8'h46 == io_in_0 ? 8'h89 : _GEN_69; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_71 = 8'h47 == io_in_0 ? 8'h87 : _GEN_70; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_72 = 8'h48 == io_in_0 ? 8'hdd : _GEN_71; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_73 = 8'h49 == io_in_0 ? 8'hd3 : _GEN_72; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_74 = 8'h4a == io_in_0 ? 8'hc1 : _GEN_73; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_75 = 8'h4b == io_in_0 ? 8'hcf : _GEN_74; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_76 = 8'h4c == io_in_0 ? 8'he5 : _GEN_75; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_77 = 8'h4d == io_in_0 ? 8'heb : _GEN_76; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_78 = 8'h4e == io_in_0 ? 8'hf9 : _GEN_77; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_79 = 8'h4f == io_in_0 ? 8'hf7 : _GEN_78; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_80 = 8'h50 == io_in_0 ? 8'h4d : _GEN_79; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_81 = 8'h51 == io_in_0 ? 8'h43 : _GEN_80; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_82 = 8'h52 == io_in_0 ? 8'h51 : _GEN_81; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_83 = 8'h53 == io_in_0 ? 8'h5f : _GEN_82; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_84 = 8'h54 == io_in_0 ? 8'h75 : _GEN_83; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_85 = 8'h55 == io_in_0 ? 8'h7b : _GEN_84; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_86 = 8'h56 == io_in_0 ? 8'h69 : _GEN_85; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_87 = 8'h57 == io_in_0 ? 8'h67 : _GEN_86; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_88 = 8'h58 == io_in_0 ? 8'h3d : _GEN_87; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_89 = 8'h59 == io_in_0 ? 8'h33 : _GEN_88; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_90 = 8'h5a == io_in_0 ? 8'h21 : _GEN_89; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_91 = 8'h5b == io_in_0 ? 8'h2f : _GEN_90; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_92 = 8'h5c == io_in_0 ? 8'h5 : _GEN_91; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_93 = 8'h5d == io_in_0 ? 8'hb : _GEN_92; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_94 = 8'h5e == io_in_0 ? 8'h19 : _GEN_93; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_95 = 8'h5f == io_in_0 ? 8'h17 : _GEN_94; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_96 = 8'h60 == io_in_0 ? 8'h76 : _GEN_95; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_97 = 8'h61 == io_in_0 ? 8'h78 : _GEN_96; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_98 = 8'h62 == io_in_0 ? 8'h6a : _GEN_97; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_99 = 8'h63 == io_in_0 ? 8'h64 : _GEN_98; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_100 = 8'h64 == io_in_0 ? 8'h4e : _GEN_99; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_101 = 8'h65 == io_in_0 ? 8'h40 : _GEN_100; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_102 = 8'h66 == io_in_0 ? 8'h52 : _GEN_101; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_103 = 8'h67 == io_in_0 ? 8'h5c : _GEN_102; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_104 = 8'h68 == io_in_0 ? 8'h6 : _GEN_103; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_105 = 8'h69 == io_in_0 ? 8'h8 : _GEN_104; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_106 = 8'h6a == io_in_0 ? 8'h1a : _GEN_105; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_107 = 8'h6b == io_in_0 ? 8'h14 : _GEN_106; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_108 = 8'h6c == io_in_0 ? 8'h3e : _GEN_107; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_109 = 8'h6d == io_in_0 ? 8'h30 : _GEN_108; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_110 = 8'h6e == io_in_0 ? 8'h22 : _GEN_109; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_111 = 8'h6f == io_in_0 ? 8'h2c : _GEN_110; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_112 = 8'h70 == io_in_0 ? 8'h96 : _GEN_111; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_113 = 8'h71 == io_in_0 ? 8'h98 : _GEN_112; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_114 = 8'h72 == io_in_0 ? 8'h8a : _GEN_113; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_115 = 8'h73 == io_in_0 ? 8'h84 : _GEN_114; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_116 = 8'h74 == io_in_0 ? 8'hae : _GEN_115; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_117 = 8'h75 == io_in_0 ? 8'ha0 : _GEN_116; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_118 = 8'h76 == io_in_0 ? 8'hb2 : _GEN_117; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_119 = 8'h77 == io_in_0 ? 8'hbc : _GEN_118; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_120 = 8'h78 == io_in_0 ? 8'he6 : _GEN_119; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_121 = 8'h79 == io_in_0 ? 8'he8 : _GEN_120; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_122 = 8'h7a == io_in_0 ? 8'hfa : _GEN_121; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_123 = 8'h7b == io_in_0 ? 8'hf4 : _GEN_122; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_124 = 8'h7c == io_in_0 ? 8'hde : _GEN_123; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_125 = 8'h7d == io_in_0 ? 8'hd0 : _GEN_124; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_126 = 8'h7e == io_in_0 ? 8'hc2 : _GEN_125; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_127 = 8'h7f == io_in_0 ? 8'hcc : _GEN_126; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_128 = 8'h80 == io_in_0 ? 8'h41 : _GEN_127; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_129 = 8'h81 == io_in_0 ? 8'h4f : _GEN_128; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_130 = 8'h82 == io_in_0 ? 8'h5d : _GEN_129; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_131 = 8'h83 == io_in_0 ? 8'h53 : _GEN_130; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_132 = 8'h84 == io_in_0 ? 8'h79 : _GEN_131; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_133 = 8'h85 == io_in_0 ? 8'h77 : _GEN_132; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_134 = 8'h86 == io_in_0 ? 8'h65 : _GEN_133; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_135 = 8'h87 == io_in_0 ? 8'h6b : _GEN_134; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_136 = 8'h88 == io_in_0 ? 8'h31 : _GEN_135; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_137 = 8'h89 == io_in_0 ? 8'h3f : _GEN_136; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_138 = 8'h8a == io_in_0 ? 8'h2d : _GEN_137; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_139 = 8'h8b == io_in_0 ? 8'h23 : _GEN_138; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_140 = 8'h8c == io_in_0 ? 8'h9 : _GEN_139; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_141 = 8'h8d == io_in_0 ? 8'h7 : _GEN_140; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_142 = 8'h8e == io_in_0 ? 8'h15 : _GEN_141; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_143 = 8'h8f == io_in_0 ? 8'h1b : _GEN_142; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_144 = 8'h90 == io_in_0 ? 8'ha1 : _GEN_143; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_145 = 8'h91 == io_in_0 ? 8'haf : _GEN_144; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_146 = 8'h92 == io_in_0 ? 8'hbd : _GEN_145; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_147 = 8'h93 == io_in_0 ? 8'hb3 : _GEN_146; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_148 = 8'h94 == io_in_0 ? 8'h99 : _GEN_147; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_149 = 8'h95 == io_in_0 ? 8'h97 : _GEN_148; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_150 = 8'h96 == io_in_0 ? 8'h85 : _GEN_149; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_151 = 8'h97 == io_in_0 ? 8'h8b : _GEN_150; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_152 = 8'h98 == io_in_0 ? 8'hd1 : _GEN_151; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_153 = 8'h99 == io_in_0 ? 8'hdf : _GEN_152; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_154 = 8'h9a == io_in_0 ? 8'hcd : _GEN_153; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_155 = 8'h9b == io_in_0 ? 8'hc3 : _GEN_154; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_156 = 8'h9c == io_in_0 ? 8'he9 : _GEN_155; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_157 = 8'h9d == io_in_0 ? 8'he7 : _GEN_156; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_158 = 8'h9e == io_in_0 ? 8'hf5 : _GEN_157; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_159 = 8'h9f == io_in_0 ? 8'hfb : _GEN_158; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_160 = 8'ha0 == io_in_0 ? 8'h9a : _GEN_159; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_161 = 8'ha1 == io_in_0 ? 8'h94 : _GEN_160; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_162 = 8'ha2 == io_in_0 ? 8'h86 : _GEN_161; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_163 = 8'ha3 == io_in_0 ? 8'h88 : _GEN_162; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_164 = 8'ha4 == io_in_0 ? 8'ha2 : _GEN_163; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_165 = 8'ha5 == io_in_0 ? 8'hac : _GEN_164; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_166 = 8'ha6 == io_in_0 ? 8'hbe : _GEN_165; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_167 = 8'ha7 == io_in_0 ? 8'hb0 : _GEN_166; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_168 = 8'ha8 == io_in_0 ? 8'hea : _GEN_167; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_169 = 8'ha9 == io_in_0 ? 8'he4 : _GEN_168; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_170 = 8'haa == io_in_0 ? 8'hf6 : _GEN_169; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_171 = 8'hab == io_in_0 ? 8'hf8 : _GEN_170; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_172 = 8'hac == io_in_0 ? 8'hd2 : _GEN_171; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_173 = 8'had == io_in_0 ? 8'hdc : _GEN_172; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_174 = 8'hae == io_in_0 ? 8'hce : _GEN_173; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_175 = 8'haf == io_in_0 ? 8'hc0 : _GEN_174; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_176 = 8'hb0 == io_in_0 ? 8'h7a : _GEN_175; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_177 = 8'hb1 == io_in_0 ? 8'h74 : _GEN_176; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_178 = 8'hb2 == io_in_0 ? 8'h66 : _GEN_177; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_179 = 8'hb3 == io_in_0 ? 8'h68 : _GEN_178; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_180 = 8'hb4 == io_in_0 ? 8'h42 : _GEN_179; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_181 = 8'hb5 == io_in_0 ? 8'h4c : _GEN_180; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_182 = 8'hb6 == io_in_0 ? 8'h5e : _GEN_181; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_183 = 8'hb7 == io_in_0 ? 8'h50 : _GEN_182; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_184 = 8'hb8 == io_in_0 ? 8'ha : _GEN_183; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_185 = 8'hb9 == io_in_0 ? 8'h4 : _GEN_184; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_186 = 8'hba == io_in_0 ? 8'h16 : _GEN_185; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_187 = 8'hbb == io_in_0 ? 8'h18 : _GEN_186; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_188 = 8'hbc == io_in_0 ? 8'h32 : _GEN_187; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_189 = 8'hbd == io_in_0 ? 8'h3c : _GEN_188; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_190 = 8'hbe == io_in_0 ? 8'h2e : _GEN_189; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_191 = 8'hbf == io_in_0 ? 8'h20 : _GEN_190; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_192 = 8'hc0 == io_in_0 ? 8'hec : _GEN_191; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_193 = 8'hc1 == io_in_0 ? 8'he2 : _GEN_192; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_194 = 8'hc2 == io_in_0 ? 8'hf0 : _GEN_193; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_195 = 8'hc3 == io_in_0 ? 8'hfe : _GEN_194; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_196 = 8'hc4 == io_in_0 ? 8'hd4 : _GEN_195; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_197 = 8'hc5 == io_in_0 ? 8'hda : _GEN_196; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_198 = 8'hc6 == io_in_0 ? 8'hc8 : _GEN_197; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_199 = 8'hc7 == io_in_0 ? 8'hc6 : _GEN_198; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_200 = 8'hc8 == io_in_0 ? 8'h9c : _GEN_199; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_201 = 8'hc9 == io_in_0 ? 8'h92 : _GEN_200; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_202 = 8'hca == io_in_0 ? 8'h80 : _GEN_201; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_203 = 8'hcb == io_in_0 ? 8'h8e : _GEN_202; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_204 = 8'hcc == io_in_0 ? 8'ha4 : _GEN_203; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_205 = 8'hcd == io_in_0 ? 8'haa : _GEN_204; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_206 = 8'hce == io_in_0 ? 8'hb8 : _GEN_205; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_207 = 8'hcf == io_in_0 ? 8'hb6 : _GEN_206; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_208 = 8'hd0 == io_in_0 ? 8'hc : _GEN_207; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_209 = 8'hd1 == io_in_0 ? 8'h2 : _GEN_208; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_210 = 8'hd2 == io_in_0 ? 8'h10 : _GEN_209; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_211 = 8'hd3 == io_in_0 ? 8'h1e : _GEN_210; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_212 = 8'hd4 == io_in_0 ? 8'h34 : _GEN_211; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_213 = 8'hd5 == io_in_0 ? 8'h3a : _GEN_212; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_214 = 8'hd6 == io_in_0 ? 8'h28 : _GEN_213; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_215 = 8'hd7 == io_in_0 ? 8'h26 : _GEN_214; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_216 = 8'hd8 == io_in_0 ? 8'h7c : _GEN_215; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_217 = 8'hd9 == io_in_0 ? 8'h72 : _GEN_216; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_218 = 8'hda == io_in_0 ? 8'h60 : _GEN_217; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_219 = 8'hdb == io_in_0 ? 8'h6e : _GEN_218; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_220 = 8'hdc == io_in_0 ? 8'h44 : _GEN_219; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_221 = 8'hdd == io_in_0 ? 8'h4a : _GEN_220; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_222 = 8'hde == io_in_0 ? 8'h58 : _GEN_221; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_223 = 8'hdf == io_in_0 ? 8'h56 : _GEN_222; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_224 = 8'he0 == io_in_0 ? 8'h37 : _GEN_223; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_225 = 8'he1 == io_in_0 ? 8'h39 : _GEN_224; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_226 = 8'he2 == io_in_0 ? 8'h2b : _GEN_225; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_227 = 8'he3 == io_in_0 ? 8'h25 : _GEN_226; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_228 = 8'he4 == io_in_0 ? 8'hf : _GEN_227; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_229 = 8'he5 == io_in_0 ? 8'h1 : _GEN_228; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_230 = 8'he6 == io_in_0 ? 8'h13 : _GEN_229; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_231 = 8'he7 == io_in_0 ? 8'h1d : _GEN_230; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_232 = 8'he8 == io_in_0 ? 8'h47 : _GEN_231; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_233 = 8'he9 == io_in_0 ? 8'h49 : _GEN_232; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_234 = 8'hea == io_in_0 ? 8'h5b : _GEN_233; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_235 = 8'heb == io_in_0 ? 8'h55 : _GEN_234; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_236 = 8'hec == io_in_0 ? 8'h7f : _GEN_235; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_237 = 8'hed == io_in_0 ? 8'h71 : _GEN_236; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_238 = 8'hee == io_in_0 ? 8'h63 : _GEN_237; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_239 = 8'hef == io_in_0 ? 8'h6d : _GEN_238; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_240 = 8'hf0 == io_in_0 ? 8'hd7 : _GEN_239; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_241 = 8'hf1 == io_in_0 ? 8'hd9 : _GEN_240; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_242 = 8'hf2 == io_in_0 ? 8'hcb : _GEN_241; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_243 = 8'hf3 == io_in_0 ? 8'hc5 : _GEN_242; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_244 = 8'hf4 == io_in_0 ? 8'hef : _GEN_243; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_245 = 8'hf5 == io_in_0 ? 8'he1 : _GEN_244; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_246 = 8'hf6 == io_in_0 ? 8'hf3 : _GEN_245; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_247 = 8'hf7 == io_in_0 ? 8'hfd : _GEN_246; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_248 = 8'hf8 == io_in_0 ? 8'ha7 : _GEN_247; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_249 = 8'hf9 == io_in_0 ? 8'ha9 : _GEN_248; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_250 = 8'hfa == io_in_0 ? 8'hbb : _GEN_249; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_251 = 8'hfb == io_in_0 ? 8'hb5 : _GEN_250; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_252 = 8'hfc == io_in_0 ? 8'h9f : _GEN_251; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_253 = 8'hfd == io_in_0 ? 8'h91 : _GEN_252; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_254 = 8'hfe == io_in_0 ? 8'h83 : _GEN_253; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_255 = 8'hff == io_in_0 ? 8'h8d : _GEN_254; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_257 = 8'h1 == io_in_1 ? 8'hb : 8'h0; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_258 = 8'h2 == io_in_1 ? 8'h16 : _GEN_257; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_259 = 8'h3 == io_in_1 ? 8'h1d : _GEN_258; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_260 = 8'h4 == io_in_1 ? 8'h2c : _GEN_259; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_261 = 8'h5 == io_in_1 ? 8'h27 : _GEN_260; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_262 = 8'h6 == io_in_1 ? 8'h3a : _GEN_261; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_263 = 8'h7 == io_in_1 ? 8'h31 : _GEN_262; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_264 = 8'h8 == io_in_1 ? 8'h58 : _GEN_263; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_265 = 8'h9 == io_in_1 ? 8'h53 : _GEN_264; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_266 = 8'ha == io_in_1 ? 8'h4e : _GEN_265; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_267 = 8'hb == io_in_1 ? 8'h45 : _GEN_266; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_268 = 8'hc == io_in_1 ? 8'h74 : _GEN_267; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_269 = 8'hd == io_in_1 ? 8'h7f : _GEN_268; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_270 = 8'he == io_in_1 ? 8'h62 : _GEN_269; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_271 = 8'hf == io_in_1 ? 8'h69 : _GEN_270; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_272 = 8'h10 == io_in_1 ? 8'hb0 : _GEN_271; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_273 = 8'h11 == io_in_1 ? 8'hbb : _GEN_272; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_274 = 8'h12 == io_in_1 ? 8'ha6 : _GEN_273; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_275 = 8'h13 == io_in_1 ? 8'had : _GEN_274; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_276 = 8'h14 == io_in_1 ? 8'h9c : _GEN_275; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_277 = 8'h15 == io_in_1 ? 8'h97 : _GEN_276; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_278 = 8'h16 == io_in_1 ? 8'h8a : _GEN_277; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_279 = 8'h17 == io_in_1 ? 8'h81 : _GEN_278; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_280 = 8'h18 == io_in_1 ? 8'he8 : _GEN_279; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_281 = 8'h19 == io_in_1 ? 8'he3 : _GEN_280; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_282 = 8'h1a == io_in_1 ? 8'hfe : _GEN_281; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_283 = 8'h1b == io_in_1 ? 8'hf5 : _GEN_282; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_284 = 8'h1c == io_in_1 ? 8'hc4 : _GEN_283; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_285 = 8'h1d == io_in_1 ? 8'hcf : _GEN_284; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_286 = 8'h1e == io_in_1 ? 8'hd2 : _GEN_285; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_287 = 8'h1f == io_in_1 ? 8'hd9 : _GEN_286; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_288 = 8'h20 == io_in_1 ? 8'h7b : _GEN_287; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_289 = 8'h21 == io_in_1 ? 8'h70 : _GEN_288; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_290 = 8'h22 == io_in_1 ? 8'h6d : _GEN_289; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_291 = 8'h23 == io_in_1 ? 8'h66 : _GEN_290; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_292 = 8'h24 == io_in_1 ? 8'h57 : _GEN_291; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_293 = 8'h25 == io_in_1 ? 8'h5c : _GEN_292; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_294 = 8'h26 == io_in_1 ? 8'h41 : _GEN_293; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_295 = 8'h27 == io_in_1 ? 8'h4a : _GEN_294; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_296 = 8'h28 == io_in_1 ? 8'h23 : _GEN_295; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_297 = 8'h29 == io_in_1 ? 8'h28 : _GEN_296; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_298 = 8'h2a == io_in_1 ? 8'h35 : _GEN_297; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_299 = 8'h2b == io_in_1 ? 8'h3e : _GEN_298; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_300 = 8'h2c == io_in_1 ? 8'hf : _GEN_299; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_301 = 8'h2d == io_in_1 ? 8'h4 : _GEN_300; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_302 = 8'h2e == io_in_1 ? 8'h19 : _GEN_301; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_303 = 8'h2f == io_in_1 ? 8'h12 : _GEN_302; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_304 = 8'h30 == io_in_1 ? 8'hcb : _GEN_303; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_305 = 8'h31 == io_in_1 ? 8'hc0 : _GEN_304; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_306 = 8'h32 == io_in_1 ? 8'hdd : _GEN_305; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_307 = 8'h33 == io_in_1 ? 8'hd6 : _GEN_306; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_308 = 8'h34 == io_in_1 ? 8'he7 : _GEN_307; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_309 = 8'h35 == io_in_1 ? 8'hec : _GEN_308; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_310 = 8'h36 == io_in_1 ? 8'hf1 : _GEN_309; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_311 = 8'h37 == io_in_1 ? 8'hfa : _GEN_310; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_312 = 8'h38 == io_in_1 ? 8'h93 : _GEN_311; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_313 = 8'h39 == io_in_1 ? 8'h98 : _GEN_312; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_314 = 8'h3a == io_in_1 ? 8'h85 : _GEN_313; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_315 = 8'h3b == io_in_1 ? 8'h8e : _GEN_314; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_316 = 8'h3c == io_in_1 ? 8'hbf : _GEN_315; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_317 = 8'h3d == io_in_1 ? 8'hb4 : _GEN_316; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_318 = 8'h3e == io_in_1 ? 8'ha9 : _GEN_317; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_319 = 8'h3f == io_in_1 ? 8'ha2 : _GEN_318; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_320 = 8'h40 == io_in_1 ? 8'hf6 : _GEN_319; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_321 = 8'h41 == io_in_1 ? 8'hfd : _GEN_320; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_322 = 8'h42 == io_in_1 ? 8'he0 : _GEN_321; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_323 = 8'h43 == io_in_1 ? 8'heb : _GEN_322; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_324 = 8'h44 == io_in_1 ? 8'hda : _GEN_323; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_325 = 8'h45 == io_in_1 ? 8'hd1 : _GEN_324; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_326 = 8'h46 == io_in_1 ? 8'hcc : _GEN_325; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_327 = 8'h47 == io_in_1 ? 8'hc7 : _GEN_326; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_328 = 8'h48 == io_in_1 ? 8'hae : _GEN_327; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_329 = 8'h49 == io_in_1 ? 8'ha5 : _GEN_328; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_330 = 8'h4a == io_in_1 ? 8'hb8 : _GEN_329; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_331 = 8'h4b == io_in_1 ? 8'hb3 : _GEN_330; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_332 = 8'h4c == io_in_1 ? 8'h82 : _GEN_331; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_333 = 8'h4d == io_in_1 ? 8'h89 : _GEN_332; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_334 = 8'h4e == io_in_1 ? 8'h94 : _GEN_333; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_335 = 8'h4f == io_in_1 ? 8'h9f : _GEN_334; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_336 = 8'h50 == io_in_1 ? 8'h46 : _GEN_335; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_337 = 8'h51 == io_in_1 ? 8'h4d : _GEN_336; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_338 = 8'h52 == io_in_1 ? 8'h50 : _GEN_337; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_339 = 8'h53 == io_in_1 ? 8'h5b : _GEN_338; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_340 = 8'h54 == io_in_1 ? 8'h6a : _GEN_339; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_341 = 8'h55 == io_in_1 ? 8'h61 : _GEN_340; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_342 = 8'h56 == io_in_1 ? 8'h7c : _GEN_341; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_343 = 8'h57 == io_in_1 ? 8'h77 : _GEN_342; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_344 = 8'h58 == io_in_1 ? 8'h1e : _GEN_343; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_345 = 8'h59 == io_in_1 ? 8'h15 : _GEN_344; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_346 = 8'h5a == io_in_1 ? 8'h8 : _GEN_345; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_347 = 8'h5b == io_in_1 ? 8'h3 : _GEN_346; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_348 = 8'h5c == io_in_1 ? 8'h32 : _GEN_347; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_349 = 8'h5d == io_in_1 ? 8'h39 : _GEN_348; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_350 = 8'h5e == io_in_1 ? 8'h24 : _GEN_349; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_351 = 8'h5f == io_in_1 ? 8'h2f : _GEN_350; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_352 = 8'h60 == io_in_1 ? 8'h8d : _GEN_351; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_353 = 8'h61 == io_in_1 ? 8'h86 : _GEN_352; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_354 = 8'h62 == io_in_1 ? 8'h9b : _GEN_353; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_355 = 8'h63 == io_in_1 ? 8'h90 : _GEN_354; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_356 = 8'h64 == io_in_1 ? 8'ha1 : _GEN_355; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_357 = 8'h65 == io_in_1 ? 8'haa : _GEN_356; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_358 = 8'h66 == io_in_1 ? 8'hb7 : _GEN_357; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_359 = 8'h67 == io_in_1 ? 8'hbc : _GEN_358; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_360 = 8'h68 == io_in_1 ? 8'hd5 : _GEN_359; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_361 = 8'h69 == io_in_1 ? 8'hde : _GEN_360; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_362 = 8'h6a == io_in_1 ? 8'hc3 : _GEN_361; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_363 = 8'h6b == io_in_1 ? 8'hc8 : _GEN_362; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_364 = 8'h6c == io_in_1 ? 8'hf9 : _GEN_363; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_365 = 8'h6d == io_in_1 ? 8'hf2 : _GEN_364; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_366 = 8'h6e == io_in_1 ? 8'hef : _GEN_365; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_367 = 8'h6f == io_in_1 ? 8'he4 : _GEN_366; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_368 = 8'h70 == io_in_1 ? 8'h3d : _GEN_367; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_369 = 8'h71 == io_in_1 ? 8'h36 : _GEN_368; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_370 = 8'h72 == io_in_1 ? 8'h2b : _GEN_369; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_371 = 8'h73 == io_in_1 ? 8'h20 : _GEN_370; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_372 = 8'h74 == io_in_1 ? 8'h11 : _GEN_371; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_373 = 8'h75 == io_in_1 ? 8'h1a : _GEN_372; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_374 = 8'h76 == io_in_1 ? 8'h7 : _GEN_373; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_375 = 8'h77 == io_in_1 ? 8'hc : _GEN_374; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_376 = 8'h78 == io_in_1 ? 8'h65 : _GEN_375; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_377 = 8'h79 == io_in_1 ? 8'h6e : _GEN_376; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_378 = 8'h7a == io_in_1 ? 8'h73 : _GEN_377; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_379 = 8'h7b == io_in_1 ? 8'h78 : _GEN_378; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_380 = 8'h7c == io_in_1 ? 8'h49 : _GEN_379; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_381 = 8'h7d == io_in_1 ? 8'h42 : _GEN_380; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_382 = 8'h7e == io_in_1 ? 8'h5f : _GEN_381; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_383 = 8'h7f == io_in_1 ? 8'h54 : _GEN_382; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_384 = 8'h80 == io_in_1 ? 8'hf7 : _GEN_383; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_385 = 8'h81 == io_in_1 ? 8'hfc : _GEN_384; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_386 = 8'h82 == io_in_1 ? 8'he1 : _GEN_385; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_387 = 8'h83 == io_in_1 ? 8'hea : _GEN_386; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_388 = 8'h84 == io_in_1 ? 8'hdb : _GEN_387; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_389 = 8'h85 == io_in_1 ? 8'hd0 : _GEN_388; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_390 = 8'h86 == io_in_1 ? 8'hcd : _GEN_389; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_391 = 8'h87 == io_in_1 ? 8'hc6 : _GEN_390; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_392 = 8'h88 == io_in_1 ? 8'haf : _GEN_391; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_393 = 8'h89 == io_in_1 ? 8'ha4 : _GEN_392; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_394 = 8'h8a == io_in_1 ? 8'hb9 : _GEN_393; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_395 = 8'h8b == io_in_1 ? 8'hb2 : _GEN_394; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_396 = 8'h8c == io_in_1 ? 8'h83 : _GEN_395; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_397 = 8'h8d == io_in_1 ? 8'h88 : _GEN_396; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_398 = 8'h8e == io_in_1 ? 8'h95 : _GEN_397; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_399 = 8'h8f == io_in_1 ? 8'h9e : _GEN_398; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_400 = 8'h90 == io_in_1 ? 8'h47 : _GEN_399; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_401 = 8'h91 == io_in_1 ? 8'h4c : _GEN_400; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_402 = 8'h92 == io_in_1 ? 8'h51 : _GEN_401; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_403 = 8'h93 == io_in_1 ? 8'h5a : _GEN_402; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_404 = 8'h94 == io_in_1 ? 8'h6b : _GEN_403; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_405 = 8'h95 == io_in_1 ? 8'h60 : _GEN_404; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_406 = 8'h96 == io_in_1 ? 8'h7d : _GEN_405; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_407 = 8'h97 == io_in_1 ? 8'h76 : _GEN_406; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_408 = 8'h98 == io_in_1 ? 8'h1f : _GEN_407; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_409 = 8'h99 == io_in_1 ? 8'h14 : _GEN_408; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_410 = 8'h9a == io_in_1 ? 8'h9 : _GEN_409; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_411 = 8'h9b == io_in_1 ? 8'h2 : _GEN_410; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_412 = 8'h9c == io_in_1 ? 8'h33 : _GEN_411; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_413 = 8'h9d == io_in_1 ? 8'h38 : _GEN_412; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_414 = 8'h9e == io_in_1 ? 8'h25 : _GEN_413; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_415 = 8'h9f == io_in_1 ? 8'h2e : _GEN_414; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_416 = 8'ha0 == io_in_1 ? 8'h8c : _GEN_415; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_417 = 8'ha1 == io_in_1 ? 8'h87 : _GEN_416; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_418 = 8'ha2 == io_in_1 ? 8'h9a : _GEN_417; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_419 = 8'ha3 == io_in_1 ? 8'h91 : _GEN_418; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_420 = 8'ha4 == io_in_1 ? 8'ha0 : _GEN_419; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_421 = 8'ha5 == io_in_1 ? 8'hab : _GEN_420; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_422 = 8'ha6 == io_in_1 ? 8'hb6 : _GEN_421; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_423 = 8'ha7 == io_in_1 ? 8'hbd : _GEN_422; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_424 = 8'ha8 == io_in_1 ? 8'hd4 : _GEN_423; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_425 = 8'ha9 == io_in_1 ? 8'hdf : _GEN_424; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_426 = 8'haa == io_in_1 ? 8'hc2 : _GEN_425; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_427 = 8'hab == io_in_1 ? 8'hc9 : _GEN_426; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_428 = 8'hac == io_in_1 ? 8'hf8 : _GEN_427; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_429 = 8'had == io_in_1 ? 8'hf3 : _GEN_428; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_430 = 8'hae == io_in_1 ? 8'hee : _GEN_429; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_431 = 8'haf == io_in_1 ? 8'he5 : _GEN_430; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_432 = 8'hb0 == io_in_1 ? 8'h3c : _GEN_431; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_433 = 8'hb1 == io_in_1 ? 8'h37 : _GEN_432; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_434 = 8'hb2 == io_in_1 ? 8'h2a : _GEN_433; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_435 = 8'hb3 == io_in_1 ? 8'h21 : _GEN_434; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_436 = 8'hb4 == io_in_1 ? 8'h10 : _GEN_435; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_437 = 8'hb5 == io_in_1 ? 8'h1b : _GEN_436; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_438 = 8'hb6 == io_in_1 ? 8'h6 : _GEN_437; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_439 = 8'hb7 == io_in_1 ? 8'hd : _GEN_438; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_440 = 8'hb8 == io_in_1 ? 8'h64 : _GEN_439; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_441 = 8'hb9 == io_in_1 ? 8'h6f : _GEN_440; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_442 = 8'hba == io_in_1 ? 8'h72 : _GEN_441; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_443 = 8'hbb == io_in_1 ? 8'h79 : _GEN_442; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_444 = 8'hbc == io_in_1 ? 8'h48 : _GEN_443; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_445 = 8'hbd == io_in_1 ? 8'h43 : _GEN_444; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_446 = 8'hbe == io_in_1 ? 8'h5e : _GEN_445; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_447 = 8'hbf == io_in_1 ? 8'h55 : _GEN_446; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_448 = 8'hc0 == io_in_1 ? 8'h1 : _GEN_447; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_449 = 8'hc1 == io_in_1 ? 8'ha : _GEN_448; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_450 = 8'hc2 == io_in_1 ? 8'h17 : _GEN_449; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_451 = 8'hc3 == io_in_1 ? 8'h1c : _GEN_450; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_452 = 8'hc4 == io_in_1 ? 8'h2d : _GEN_451; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_453 = 8'hc5 == io_in_1 ? 8'h26 : _GEN_452; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_454 = 8'hc6 == io_in_1 ? 8'h3b : _GEN_453; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_455 = 8'hc7 == io_in_1 ? 8'h30 : _GEN_454; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_456 = 8'hc8 == io_in_1 ? 8'h59 : _GEN_455; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_457 = 8'hc9 == io_in_1 ? 8'h52 : _GEN_456; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_458 = 8'hca == io_in_1 ? 8'h4f : _GEN_457; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_459 = 8'hcb == io_in_1 ? 8'h44 : _GEN_458; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_460 = 8'hcc == io_in_1 ? 8'h75 : _GEN_459; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_461 = 8'hcd == io_in_1 ? 8'h7e : _GEN_460; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_462 = 8'hce == io_in_1 ? 8'h63 : _GEN_461; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_463 = 8'hcf == io_in_1 ? 8'h68 : _GEN_462; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_464 = 8'hd0 == io_in_1 ? 8'hb1 : _GEN_463; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_465 = 8'hd1 == io_in_1 ? 8'hba : _GEN_464; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_466 = 8'hd2 == io_in_1 ? 8'ha7 : _GEN_465; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_467 = 8'hd3 == io_in_1 ? 8'hac : _GEN_466; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_468 = 8'hd4 == io_in_1 ? 8'h9d : _GEN_467; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_469 = 8'hd5 == io_in_1 ? 8'h96 : _GEN_468; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_470 = 8'hd6 == io_in_1 ? 8'h8b : _GEN_469; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_471 = 8'hd7 == io_in_1 ? 8'h80 : _GEN_470; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_472 = 8'hd8 == io_in_1 ? 8'he9 : _GEN_471; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_473 = 8'hd9 == io_in_1 ? 8'he2 : _GEN_472; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_474 = 8'hda == io_in_1 ? 8'hff : _GEN_473; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_475 = 8'hdb == io_in_1 ? 8'hf4 : _GEN_474; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_476 = 8'hdc == io_in_1 ? 8'hc5 : _GEN_475; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_477 = 8'hdd == io_in_1 ? 8'hce : _GEN_476; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_478 = 8'hde == io_in_1 ? 8'hd3 : _GEN_477; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_479 = 8'hdf == io_in_1 ? 8'hd8 : _GEN_478; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_480 = 8'he0 == io_in_1 ? 8'h7a : _GEN_479; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_481 = 8'he1 == io_in_1 ? 8'h71 : _GEN_480; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_482 = 8'he2 == io_in_1 ? 8'h6c : _GEN_481; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_483 = 8'he3 == io_in_1 ? 8'h67 : _GEN_482; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_484 = 8'he4 == io_in_1 ? 8'h56 : _GEN_483; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_485 = 8'he5 == io_in_1 ? 8'h5d : _GEN_484; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_486 = 8'he6 == io_in_1 ? 8'h40 : _GEN_485; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_487 = 8'he7 == io_in_1 ? 8'h4b : _GEN_486; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_488 = 8'he8 == io_in_1 ? 8'h22 : _GEN_487; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_489 = 8'he9 == io_in_1 ? 8'h29 : _GEN_488; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_490 = 8'hea == io_in_1 ? 8'h34 : _GEN_489; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_491 = 8'heb == io_in_1 ? 8'h3f : _GEN_490; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_492 = 8'hec == io_in_1 ? 8'he : _GEN_491; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_493 = 8'hed == io_in_1 ? 8'h5 : _GEN_492; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_494 = 8'hee == io_in_1 ? 8'h18 : _GEN_493; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_495 = 8'hef == io_in_1 ? 8'h13 : _GEN_494; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_496 = 8'hf0 == io_in_1 ? 8'hca : _GEN_495; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_497 = 8'hf1 == io_in_1 ? 8'hc1 : _GEN_496; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_498 = 8'hf2 == io_in_1 ? 8'hdc : _GEN_497; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_499 = 8'hf3 == io_in_1 ? 8'hd7 : _GEN_498; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_500 = 8'hf4 == io_in_1 ? 8'he6 : _GEN_499; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_501 = 8'hf5 == io_in_1 ? 8'hed : _GEN_500; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_502 = 8'hf6 == io_in_1 ? 8'hf0 : _GEN_501; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_503 = 8'hf7 == io_in_1 ? 8'hfb : _GEN_502; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_504 = 8'hf8 == io_in_1 ? 8'h92 : _GEN_503; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_505 = 8'hf9 == io_in_1 ? 8'h99 : _GEN_504; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_506 = 8'hfa == io_in_1 ? 8'h84 : _GEN_505; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_507 = 8'hfb == io_in_1 ? 8'h8f : _GEN_506; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_508 = 8'hfc == io_in_1 ? 8'hbe : _GEN_507; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_509 = 8'hfd == io_in_1 ? 8'hb5 : _GEN_508; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_510 = 8'hfe == io_in_1 ? 8'ha8 : _GEN_509; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_511 = 8'hff == io_in_1 ? 8'ha3 : _GEN_510; // @[AES_PipelinedElasticBuffer.scala 591:32 AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _T = _GEN_255 ^ _GEN_511; // @[AES_PipelinedElasticBuffer.scala 591:32]
  wire [7:0] _GEN_513 = 8'h1 == io_in_2 ? 8'hd : 8'h0; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_514 = 8'h2 == io_in_2 ? 8'h1a : _GEN_513; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_515 = 8'h3 == io_in_2 ? 8'h17 : _GEN_514; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_516 = 8'h4 == io_in_2 ? 8'h34 : _GEN_515; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_517 = 8'h5 == io_in_2 ? 8'h39 : _GEN_516; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_518 = 8'h6 == io_in_2 ? 8'h2e : _GEN_517; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_519 = 8'h7 == io_in_2 ? 8'h23 : _GEN_518; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_520 = 8'h8 == io_in_2 ? 8'h68 : _GEN_519; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_521 = 8'h9 == io_in_2 ? 8'h65 : _GEN_520; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_522 = 8'ha == io_in_2 ? 8'h72 : _GEN_521; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_523 = 8'hb == io_in_2 ? 8'h7f : _GEN_522; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_524 = 8'hc == io_in_2 ? 8'h5c : _GEN_523; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_525 = 8'hd == io_in_2 ? 8'h51 : _GEN_524; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_526 = 8'he == io_in_2 ? 8'h46 : _GEN_525; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_527 = 8'hf == io_in_2 ? 8'h4b : _GEN_526; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_528 = 8'h10 == io_in_2 ? 8'hd0 : _GEN_527; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_529 = 8'h11 == io_in_2 ? 8'hdd : _GEN_528; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_530 = 8'h12 == io_in_2 ? 8'hca : _GEN_529; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_531 = 8'h13 == io_in_2 ? 8'hc7 : _GEN_530; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_532 = 8'h14 == io_in_2 ? 8'he4 : _GEN_531; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_533 = 8'h15 == io_in_2 ? 8'he9 : _GEN_532; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_534 = 8'h16 == io_in_2 ? 8'hfe : _GEN_533; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_535 = 8'h17 == io_in_2 ? 8'hf3 : _GEN_534; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_536 = 8'h18 == io_in_2 ? 8'hb8 : _GEN_535; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_537 = 8'h19 == io_in_2 ? 8'hb5 : _GEN_536; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_538 = 8'h1a == io_in_2 ? 8'ha2 : _GEN_537; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_539 = 8'h1b == io_in_2 ? 8'haf : _GEN_538; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_540 = 8'h1c == io_in_2 ? 8'h8c : _GEN_539; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_541 = 8'h1d == io_in_2 ? 8'h81 : _GEN_540; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_542 = 8'h1e == io_in_2 ? 8'h96 : _GEN_541; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_543 = 8'h1f == io_in_2 ? 8'h9b : _GEN_542; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_544 = 8'h20 == io_in_2 ? 8'hbb : _GEN_543; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_545 = 8'h21 == io_in_2 ? 8'hb6 : _GEN_544; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_546 = 8'h22 == io_in_2 ? 8'ha1 : _GEN_545; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_547 = 8'h23 == io_in_2 ? 8'hac : _GEN_546; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_548 = 8'h24 == io_in_2 ? 8'h8f : _GEN_547; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_549 = 8'h25 == io_in_2 ? 8'h82 : _GEN_548; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_550 = 8'h26 == io_in_2 ? 8'h95 : _GEN_549; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_551 = 8'h27 == io_in_2 ? 8'h98 : _GEN_550; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_552 = 8'h28 == io_in_2 ? 8'hd3 : _GEN_551; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_553 = 8'h29 == io_in_2 ? 8'hde : _GEN_552; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_554 = 8'h2a == io_in_2 ? 8'hc9 : _GEN_553; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_555 = 8'h2b == io_in_2 ? 8'hc4 : _GEN_554; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_556 = 8'h2c == io_in_2 ? 8'he7 : _GEN_555; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_557 = 8'h2d == io_in_2 ? 8'hea : _GEN_556; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_558 = 8'h2e == io_in_2 ? 8'hfd : _GEN_557; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_559 = 8'h2f == io_in_2 ? 8'hf0 : _GEN_558; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_560 = 8'h30 == io_in_2 ? 8'h6b : _GEN_559; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_561 = 8'h31 == io_in_2 ? 8'h66 : _GEN_560; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_562 = 8'h32 == io_in_2 ? 8'h71 : _GEN_561; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_563 = 8'h33 == io_in_2 ? 8'h7c : _GEN_562; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_564 = 8'h34 == io_in_2 ? 8'h5f : _GEN_563; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_565 = 8'h35 == io_in_2 ? 8'h52 : _GEN_564; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_566 = 8'h36 == io_in_2 ? 8'h45 : _GEN_565; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_567 = 8'h37 == io_in_2 ? 8'h48 : _GEN_566; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_568 = 8'h38 == io_in_2 ? 8'h3 : _GEN_567; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_569 = 8'h39 == io_in_2 ? 8'he : _GEN_568; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_570 = 8'h3a == io_in_2 ? 8'h19 : _GEN_569; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_571 = 8'h3b == io_in_2 ? 8'h14 : _GEN_570; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_572 = 8'h3c == io_in_2 ? 8'h37 : _GEN_571; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_573 = 8'h3d == io_in_2 ? 8'h3a : _GEN_572; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_574 = 8'h3e == io_in_2 ? 8'h2d : _GEN_573; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_575 = 8'h3f == io_in_2 ? 8'h20 : _GEN_574; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_576 = 8'h40 == io_in_2 ? 8'h6d : _GEN_575; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_577 = 8'h41 == io_in_2 ? 8'h60 : _GEN_576; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_578 = 8'h42 == io_in_2 ? 8'h77 : _GEN_577; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_579 = 8'h43 == io_in_2 ? 8'h7a : _GEN_578; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_580 = 8'h44 == io_in_2 ? 8'h59 : _GEN_579; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_581 = 8'h45 == io_in_2 ? 8'h54 : _GEN_580; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_582 = 8'h46 == io_in_2 ? 8'h43 : _GEN_581; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_583 = 8'h47 == io_in_2 ? 8'h4e : _GEN_582; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_584 = 8'h48 == io_in_2 ? 8'h5 : _GEN_583; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_585 = 8'h49 == io_in_2 ? 8'h8 : _GEN_584; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_586 = 8'h4a == io_in_2 ? 8'h1f : _GEN_585; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_587 = 8'h4b == io_in_2 ? 8'h12 : _GEN_586; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_588 = 8'h4c == io_in_2 ? 8'h31 : _GEN_587; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_589 = 8'h4d == io_in_2 ? 8'h3c : _GEN_588; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_590 = 8'h4e == io_in_2 ? 8'h2b : _GEN_589; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_591 = 8'h4f == io_in_2 ? 8'h26 : _GEN_590; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_592 = 8'h50 == io_in_2 ? 8'hbd : _GEN_591; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_593 = 8'h51 == io_in_2 ? 8'hb0 : _GEN_592; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_594 = 8'h52 == io_in_2 ? 8'ha7 : _GEN_593; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_595 = 8'h53 == io_in_2 ? 8'haa : _GEN_594; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_596 = 8'h54 == io_in_2 ? 8'h89 : _GEN_595; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_597 = 8'h55 == io_in_2 ? 8'h84 : _GEN_596; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_598 = 8'h56 == io_in_2 ? 8'h93 : _GEN_597; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_599 = 8'h57 == io_in_2 ? 8'h9e : _GEN_598; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_600 = 8'h58 == io_in_2 ? 8'hd5 : _GEN_599; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_601 = 8'h59 == io_in_2 ? 8'hd8 : _GEN_600; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_602 = 8'h5a == io_in_2 ? 8'hcf : _GEN_601; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_603 = 8'h5b == io_in_2 ? 8'hc2 : _GEN_602; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_604 = 8'h5c == io_in_2 ? 8'he1 : _GEN_603; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_605 = 8'h5d == io_in_2 ? 8'hec : _GEN_604; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_606 = 8'h5e == io_in_2 ? 8'hfb : _GEN_605; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_607 = 8'h5f == io_in_2 ? 8'hf6 : _GEN_606; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_608 = 8'h60 == io_in_2 ? 8'hd6 : _GEN_607; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_609 = 8'h61 == io_in_2 ? 8'hdb : _GEN_608; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_610 = 8'h62 == io_in_2 ? 8'hcc : _GEN_609; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_611 = 8'h63 == io_in_2 ? 8'hc1 : _GEN_610; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_612 = 8'h64 == io_in_2 ? 8'he2 : _GEN_611; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_613 = 8'h65 == io_in_2 ? 8'hef : _GEN_612; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_614 = 8'h66 == io_in_2 ? 8'hf8 : _GEN_613; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_615 = 8'h67 == io_in_2 ? 8'hf5 : _GEN_614; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_616 = 8'h68 == io_in_2 ? 8'hbe : _GEN_615; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_617 = 8'h69 == io_in_2 ? 8'hb3 : _GEN_616; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_618 = 8'h6a == io_in_2 ? 8'ha4 : _GEN_617; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_619 = 8'h6b == io_in_2 ? 8'ha9 : _GEN_618; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_620 = 8'h6c == io_in_2 ? 8'h8a : _GEN_619; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_621 = 8'h6d == io_in_2 ? 8'h87 : _GEN_620; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_622 = 8'h6e == io_in_2 ? 8'h90 : _GEN_621; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_623 = 8'h6f == io_in_2 ? 8'h9d : _GEN_622; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_624 = 8'h70 == io_in_2 ? 8'h6 : _GEN_623; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_625 = 8'h71 == io_in_2 ? 8'hb : _GEN_624; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_626 = 8'h72 == io_in_2 ? 8'h1c : _GEN_625; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_627 = 8'h73 == io_in_2 ? 8'h11 : _GEN_626; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_628 = 8'h74 == io_in_2 ? 8'h32 : _GEN_627; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_629 = 8'h75 == io_in_2 ? 8'h3f : _GEN_628; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_630 = 8'h76 == io_in_2 ? 8'h28 : _GEN_629; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_631 = 8'h77 == io_in_2 ? 8'h25 : _GEN_630; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_632 = 8'h78 == io_in_2 ? 8'h6e : _GEN_631; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_633 = 8'h79 == io_in_2 ? 8'h63 : _GEN_632; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_634 = 8'h7a == io_in_2 ? 8'h74 : _GEN_633; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_635 = 8'h7b == io_in_2 ? 8'h79 : _GEN_634; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_636 = 8'h7c == io_in_2 ? 8'h5a : _GEN_635; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_637 = 8'h7d == io_in_2 ? 8'h57 : _GEN_636; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_638 = 8'h7e == io_in_2 ? 8'h40 : _GEN_637; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_639 = 8'h7f == io_in_2 ? 8'h4d : _GEN_638; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_640 = 8'h80 == io_in_2 ? 8'hda : _GEN_639; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_641 = 8'h81 == io_in_2 ? 8'hd7 : _GEN_640; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_642 = 8'h82 == io_in_2 ? 8'hc0 : _GEN_641; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_643 = 8'h83 == io_in_2 ? 8'hcd : _GEN_642; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_644 = 8'h84 == io_in_2 ? 8'hee : _GEN_643; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_645 = 8'h85 == io_in_2 ? 8'he3 : _GEN_644; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_646 = 8'h86 == io_in_2 ? 8'hf4 : _GEN_645; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_647 = 8'h87 == io_in_2 ? 8'hf9 : _GEN_646; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_648 = 8'h88 == io_in_2 ? 8'hb2 : _GEN_647; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_649 = 8'h89 == io_in_2 ? 8'hbf : _GEN_648; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_650 = 8'h8a == io_in_2 ? 8'ha8 : _GEN_649; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_651 = 8'h8b == io_in_2 ? 8'ha5 : _GEN_650; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_652 = 8'h8c == io_in_2 ? 8'h86 : _GEN_651; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_653 = 8'h8d == io_in_2 ? 8'h8b : _GEN_652; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_654 = 8'h8e == io_in_2 ? 8'h9c : _GEN_653; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_655 = 8'h8f == io_in_2 ? 8'h91 : _GEN_654; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_656 = 8'h90 == io_in_2 ? 8'ha : _GEN_655; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_657 = 8'h91 == io_in_2 ? 8'h7 : _GEN_656; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_658 = 8'h92 == io_in_2 ? 8'h10 : _GEN_657; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_659 = 8'h93 == io_in_2 ? 8'h1d : _GEN_658; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_660 = 8'h94 == io_in_2 ? 8'h3e : _GEN_659; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_661 = 8'h95 == io_in_2 ? 8'h33 : _GEN_660; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_662 = 8'h96 == io_in_2 ? 8'h24 : _GEN_661; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_663 = 8'h97 == io_in_2 ? 8'h29 : _GEN_662; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_664 = 8'h98 == io_in_2 ? 8'h62 : _GEN_663; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_665 = 8'h99 == io_in_2 ? 8'h6f : _GEN_664; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_666 = 8'h9a == io_in_2 ? 8'h78 : _GEN_665; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_667 = 8'h9b == io_in_2 ? 8'h75 : _GEN_666; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_668 = 8'h9c == io_in_2 ? 8'h56 : _GEN_667; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_669 = 8'h9d == io_in_2 ? 8'h5b : _GEN_668; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_670 = 8'h9e == io_in_2 ? 8'h4c : _GEN_669; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_671 = 8'h9f == io_in_2 ? 8'h41 : _GEN_670; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_672 = 8'ha0 == io_in_2 ? 8'h61 : _GEN_671; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_673 = 8'ha1 == io_in_2 ? 8'h6c : _GEN_672; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_674 = 8'ha2 == io_in_2 ? 8'h7b : _GEN_673; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_675 = 8'ha3 == io_in_2 ? 8'h76 : _GEN_674; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_676 = 8'ha4 == io_in_2 ? 8'h55 : _GEN_675; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_677 = 8'ha5 == io_in_2 ? 8'h58 : _GEN_676; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_678 = 8'ha6 == io_in_2 ? 8'h4f : _GEN_677; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_679 = 8'ha7 == io_in_2 ? 8'h42 : _GEN_678; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_680 = 8'ha8 == io_in_2 ? 8'h9 : _GEN_679; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_681 = 8'ha9 == io_in_2 ? 8'h4 : _GEN_680; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_682 = 8'haa == io_in_2 ? 8'h13 : _GEN_681; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_683 = 8'hab == io_in_2 ? 8'h1e : _GEN_682; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_684 = 8'hac == io_in_2 ? 8'h3d : _GEN_683; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_685 = 8'had == io_in_2 ? 8'h30 : _GEN_684; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_686 = 8'hae == io_in_2 ? 8'h27 : _GEN_685; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_687 = 8'haf == io_in_2 ? 8'h2a : _GEN_686; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_688 = 8'hb0 == io_in_2 ? 8'hb1 : _GEN_687; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_689 = 8'hb1 == io_in_2 ? 8'hbc : _GEN_688; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_690 = 8'hb2 == io_in_2 ? 8'hab : _GEN_689; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_691 = 8'hb3 == io_in_2 ? 8'ha6 : _GEN_690; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_692 = 8'hb4 == io_in_2 ? 8'h85 : _GEN_691; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_693 = 8'hb5 == io_in_2 ? 8'h88 : _GEN_692; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_694 = 8'hb6 == io_in_2 ? 8'h9f : _GEN_693; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_695 = 8'hb7 == io_in_2 ? 8'h92 : _GEN_694; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_696 = 8'hb8 == io_in_2 ? 8'hd9 : _GEN_695; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_697 = 8'hb9 == io_in_2 ? 8'hd4 : _GEN_696; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_698 = 8'hba == io_in_2 ? 8'hc3 : _GEN_697; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_699 = 8'hbb == io_in_2 ? 8'hce : _GEN_698; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_700 = 8'hbc == io_in_2 ? 8'hed : _GEN_699; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_701 = 8'hbd == io_in_2 ? 8'he0 : _GEN_700; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_702 = 8'hbe == io_in_2 ? 8'hf7 : _GEN_701; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_703 = 8'hbf == io_in_2 ? 8'hfa : _GEN_702; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_704 = 8'hc0 == io_in_2 ? 8'hb7 : _GEN_703; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_705 = 8'hc1 == io_in_2 ? 8'hba : _GEN_704; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_706 = 8'hc2 == io_in_2 ? 8'had : _GEN_705; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_707 = 8'hc3 == io_in_2 ? 8'ha0 : _GEN_706; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_708 = 8'hc4 == io_in_2 ? 8'h83 : _GEN_707; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_709 = 8'hc5 == io_in_2 ? 8'h8e : _GEN_708; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_710 = 8'hc6 == io_in_2 ? 8'h99 : _GEN_709; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_711 = 8'hc7 == io_in_2 ? 8'h94 : _GEN_710; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_712 = 8'hc8 == io_in_2 ? 8'hdf : _GEN_711; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_713 = 8'hc9 == io_in_2 ? 8'hd2 : _GEN_712; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_714 = 8'hca == io_in_2 ? 8'hc5 : _GEN_713; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_715 = 8'hcb == io_in_2 ? 8'hc8 : _GEN_714; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_716 = 8'hcc == io_in_2 ? 8'heb : _GEN_715; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_717 = 8'hcd == io_in_2 ? 8'he6 : _GEN_716; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_718 = 8'hce == io_in_2 ? 8'hf1 : _GEN_717; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_719 = 8'hcf == io_in_2 ? 8'hfc : _GEN_718; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_720 = 8'hd0 == io_in_2 ? 8'h67 : _GEN_719; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_721 = 8'hd1 == io_in_2 ? 8'h6a : _GEN_720; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_722 = 8'hd2 == io_in_2 ? 8'h7d : _GEN_721; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_723 = 8'hd3 == io_in_2 ? 8'h70 : _GEN_722; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_724 = 8'hd4 == io_in_2 ? 8'h53 : _GEN_723; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_725 = 8'hd5 == io_in_2 ? 8'h5e : _GEN_724; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_726 = 8'hd6 == io_in_2 ? 8'h49 : _GEN_725; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_727 = 8'hd7 == io_in_2 ? 8'h44 : _GEN_726; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_728 = 8'hd8 == io_in_2 ? 8'hf : _GEN_727; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_729 = 8'hd9 == io_in_2 ? 8'h2 : _GEN_728; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_730 = 8'hda == io_in_2 ? 8'h15 : _GEN_729; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_731 = 8'hdb == io_in_2 ? 8'h18 : _GEN_730; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_732 = 8'hdc == io_in_2 ? 8'h3b : _GEN_731; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_733 = 8'hdd == io_in_2 ? 8'h36 : _GEN_732; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_734 = 8'hde == io_in_2 ? 8'h21 : _GEN_733; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_735 = 8'hdf == io_in_2 ? 8'h2c : _GEN_734; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_736 = 8'he0 == io_in_2 ? 8'hc : _GEN_735; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_737 = 8'he1 == io_in_2 ? 8'h1 : _GEN_736; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_738 = 8'he2 == io_in_2 ? 8'h16 : _GEN_737; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_739 = 8'he3 == io_in_2 ? 8'h1b : _GEN_738; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_740 = 8'he4 == io_in_2 ? 8'h38 : _GEN_739; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_741 = 8'he5 == io_in_2 ? 8'h35 : _GEN_740; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_742 = 8'he6 == io_in_2 ? 8'h22 : _GEN_741; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_743 = 8'he7 == io_in_2 ? 8'h2f : _GEN_742; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_744 = 8'he8 == io_in_2 ? 8'h64 : _GEN_743; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_745 = 8'he9 == io_in_2 ? 8'h69 : _GEN_744; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_746 = 8'hea == io_in_2 ? 8'h7e : _GEN_745; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_747 = 8'heb == io_in_2 ? 8'h73 : _GEN_746; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_748 = 8'hec == io_in_2 ? 8'h50 : _GEN_747; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_749 = 8'hed == io_in_2 ? 8'h5d : _GEN_748; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_750 = 8'hee == io_in_2 ? 8'h4a : _GEN_749; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_751 = 8'hef == io_in_2 ? 8'h47 : _GEN_750; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_752 = 8'hf0 == io_in_2 ? 8'hdc : _GEN_751; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_753 = 8'hf1 == io_in_2 ? 8'hd1 : _GEN_752; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_754 = 8'hf2 == io_in_2 ? 8'hc6 : _GEN_753; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_755 = 8'hf3 == io_in_2 ? 8'hcb : _GEN_754; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_756 = 8'hf4 == io_in_2 ? 8'he8 : _GEN_755; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_757 = 8'hf5 == io_in_2 ? 8'he5 : _GEN_756; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_758 = 8'hf6 == io_in_2 ? 8'hf2 : _GEN_757; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_759 = 8'hf7 == io_in_2 ? 8'hff : _GEN_758; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_760 = 8'hf8 == io_in_2 ? 8'hb4 : _GEN_759; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_761 = 8'hf9 == io_in_2 ? 8'hb9 : _GEN_760; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_762 = 8'hfa == io_in_2 ? 8'hae : _GEN_761; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_763 = 8'hfb == io_in_2 ? 8'ha3 : _GEN_762; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_764 = 8'hfc == io_in_2 ? 8'h80 : _GEN_763; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_765 = 8'hfd == io_in_2 ? 8'h8d : _GEN_764; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_766 = 8'hfe == io_in_2 ? 8'h9a : _GEN_765; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_767 = 8'hff == io_in_2 ? 8'h97 : _GEN_766; // @[AES_PipelinedElasticBuffer.scala 591:50 AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _T_1 = _T ^ _GEN_767; // @[AES_PipelinedElasticBuffer.scala 591:50]
  wire [7:0] _GEN_769 = 8'h1 == io_in_3 ? 8'h9 : 8'h0; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_770 = 8'h2 == io_in_3 ? 8'h12 : _GEN_769; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_771 = 8'h3 == io_in_3 ? 8'h1b : _GEN_770; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_772 = 8'h4 == io_in_3 ? 8'h24 : _GEN_771; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_773 = 8'h5 == io_in_3 ? 8'h2d : _GEN_772; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_774 = 8'h6 == io_in_3 ? 8'h36 : _GEN_773; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_775 = 8'h7 == io_in_3 ? 8'h3f : _GEN_774; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_776 = 8'h8 == io_in_3 ? 8'h48 : _GEN_775; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_777 = 8'h9 == io_in_3 ? 8'h41 : _GEN_776; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_778 = 8'ha == io_in_3 ? 8'h5a : _GEN_777; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_779 = 8'hb == io_in_3 ? 8'h53 : _GEN_778; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_780 = 8'hc == io_in_3 ? 8'h6c : _GEN_779; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_781 = 8'hd == io_in_3 ? 8'h65 : _GEN_780; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_782 = 8'he == io_in_3 ? 8'h7e : _GEN_781; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_783 = 8'hf == io_in_3 ? 8'h77 : _GEN_782; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_784 = 8'h10 == io_in_3 ? 8'h90 : _GEN_783; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_785 = 8'h11 == io_in_3 ? 8'h99 : _GEN_784; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_786 = 8'h12 == io_in_3 ? 8'h82 : _GEN_785; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_787 = 8'h13 == io_in_3 ? 8'h8b : _GEN_786; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_788 = 8'h14 == io_in_3 ? 8'hb4 : _GEN_787; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_789 = 8'h15 == io_in_3 ? 8'hbd : _GEN_788; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_790 = 8'h16 == io_in_3 ? 8'ha6 : _GEN_789; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_791 = 8'h17 == io_in_3 ? 8'haf : _GEN_790; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_792 = 8'h18 == io_in_3 ? 8'hd8 : _GEN_791; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_793 = 8'h19 == io_in_3 ? 8'hd1 : _GEN_792; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_794 = 8'h1a == io_in_3 ? 8'hca : _GEN_793; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_795 = 8'h1b == io_in_3 ? 8'hc3 : _GEN_794; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_796 = 8'h1c == io_in_3 ? 8'hfc : _GEN_795; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_797 = 8'h1d == io_in_3 ? 8'hf5 : _GEN_796; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_798 = 8'h1e == io_in_3 ? 8'hee : _GEN_797; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_799 = 8'h1f == io_in_3 ? 8'he7 : _GEN_798; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_800 = 8'h20 == io_in_3 ? 8'h3b : _GEN_799; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_801 = 8'h21 == io_in_3 ? 8'h32 : _GEN_800; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_802 = 8'h22 == io_in_3 ? 8'h29 : _GEN_801; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_803 = 8'h23 == io_in_3 ? 8'h20 : _GEN_802; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_804 = 8'h24 == io_in_3 ? 8'h1f : _GEN_803; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_805 = 8'h25 == io_in_3 ? 8'h16 : _GEN_804; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_806 = 8'h26 == io_in_3 ? 8'hd : _GEN_805; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_807 = 8'h27 == io_in_3 ? 8'h4 : _GEN_806; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_808 = 8'h28 == io_in_3 ? 8'h73 : _GEN_807; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_809 = 8'h29 == io_in_3 ? 8'h7a : _GEN_808; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_810 = 8'h2a == io_in_3 ? 8'h61 : _GEN_809; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_811 = 8'h2b == io_in_3 ? 8'h68 : _GEN_810; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_812 = 8'h2c == io_in_3 ? 8'h57 : _GEN_811; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_813 = 8'h2d == io_in_3 ? 8'h5e : _GEN_812; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_814 = 8'h2e == io_in_3 ? 8'h45 : _GEN_813; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_815 = 8'h2f == io_in_3 ? 8'h4c : _GEN_814; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_816 = 8'h30 == io_in_3 ? 8'hab : _GEN_815; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_817 = 8'h31 == io_in_3 ? 8'ha2 : _GEN_816; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_818 = 8'h32 == io_in_3 ? 8'hb9 : _GEN_817; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_819 = 8'h33 == io_in_3 ? 8'hb0 : _GEN_818; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_820 = 8'h34 == io_in_3 ? 8'h8f : _GEN_819; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_821 = 8'h35 == io_in_3 ? 8'h86 : _GEN_820; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_822 = 8'h36 == io_in_3 ? 8'h9d : _GEN_821; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_823 = 8'h37 == io_in_3 ? 8'h94 : _GEN_822; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_824 = 8'h38 == io_in_3 ? 8'he3 : _GEN_823; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_825 = 8'h39 == io_in_3 ? 8'hea : _GEN_824; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_826 = 8'h3a == io_in_3 ? 8'hf1 : _GEN_825; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_827 = 8'h3b == io_in_3 ? 8'hf8 : _GEN_826; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_828 = 8'h3c == io_in_3 ? 8'hc7 : _GEN_827; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_829 = 8'h3d == io_in_3 ? 8'hce : _GEN_828; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_830 = 8'h3e == io_in_3 ? 8'hd5 : _GEN_829; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_831 = 8'h3f == io_in_3 ? 8'hdc : _GEN_830; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_832 = 8'h40 == io_in_3 ? 8'h76 : _GEN_831; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_833 = 8'h41 == io_in_3 ? 8'h7f : _GEN_832; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_834 = 8'h42 == io_in_3 ? 8'h64 : _GEN_833; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_835 = 8'h43 == io_in_3 ? 8'h6d : _GEN_834; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_836 = 8'h44 == io_in_3 ? 8'h52 : _GEN_835; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_837 = 8'h45 == io_in_3 ? 8'h5b : _GEN_836; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_838 = 8'h46 == io_in_3 ? 8'h40 : _GEN_837; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_839 = 8'h47 == io_in_3 ? 8'h49 : _GEN_838; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_840 = 8'h48 == io_in_3 ? 8'h3e : _GEN_839; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_841 = 8'h49 == io_in_3 ? 8'h37 : _GEN_840; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_842 = 8'h4a == io_in_3 ? 8'h2c : _GEN_841; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_843 = 8'h4b == io_in_3 ? 8'h25 : _GEN_842; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_844 = 8'h4c == io_in_3 ? 8'h1a : _GEN_843; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_845 = 8'h4d == io_in_3 ? 8'h13 : _GEN_844; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_846 = 8'h4e == io_in_3 ? 8'h8 : _GEN_845; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_847 = 8'h4f == io_in_3 ? 8'h1 : _GEN_846; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_848 = 8'h50 == io_in_3 ? 8'he6 : _GEN_847; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_849 = 8'h51 == io_in_3 ? 8'hef : _GEN_848; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_850 = 8'h52 == io_in_3 ? 8'hf4 : _GEN_849; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_851 = 8'h53 == io_in_3 ? 8'hfd : _GEN_850; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_852 = 8'h54 == io_in_3 ? 8'hc2 : _GEN_851; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_853 = 8'h55 == io_in_3 ? 8'hcb : _GEN_852; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_854 = 8'h56 == io_in_3 ? 8'hd0 : _GEN_853; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_855 = 8'h57 == io_in_3 ? 8'hd9 : _GEN_854; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_856 = 8'h58 == io_in_3 ? 8'hae : _GEN_855; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_857 = 8'h59 == io_in_3 ? 8'ha7 : _GEN_856; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_858 = 8'h5a == io_in_3 ? 8'hbc : _GEN_857; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_859 = 8'h5b == io_in_3 ? 8'hb5 : _GEN_858; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_860 = 8'h5c == io_in_3 ? 8'h8a : _GEN_859; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_861 = 8'h5d == io_in_3 ? 8'h83 : _GEN_860; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_862 = 8'h5e == io_in_3 ? 8'h98 : _GEN_861; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_863 = 8'h5f == io_in_3 ? 8'h91 : _GEN_862; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_864 = 8'h60 == io_in_3 ? 8'h4d : _GEN_863; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_865 = 8'h61 == io_in_3 ? 8'h44 : _GEN_864; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_866 = 8'h62 == io_in_3 ? 8'h5f : _GEN_865; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_867 = 8'h63 == io_in_3 ? 8'h56 : _GEN_866; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_868 = 8'h64 == io_in_3 ? 8'h69 : _GEN_867; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_869 = 8'h65 == io_in_3 ? 8'h60 : _GEN_868; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_870 = 8'h66 == io_in_3 ? 8'h7b : _GEN_869; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_871 = 8'h67 == io_in_3 ? 8'h72 : _GEN_870; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_872 = 8'h68 == io_in_3 ? 8'h5 : _GEN_871; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_873 = 8'h69 == io_in_3 ? 8'hc : _GEN_872; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_874 = 8'h6a == io_in_3 ? 8'h17 : _GEN_873; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_875 = 8'h6b == io_in_3 ? 8'h1e : _GEN_874; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_876 = 8'h6c == io_in_3 ? 8'h21 : _GEN_875; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_877 = 8'h6d == io_in_3 ? 8'h28 : _GEN_876; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_878 = 8'h6e == io_in_3 ? 8'h33 : _GEN_877; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_879 = 8'h6f == io_in_3 ? 8'h3a : _GEN_878; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_880 = 8'h70 == io_in_3 ? 8'hdd : _GEN_879; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_881 = 8'h71 == io_in_3 ? 8'hd4 : _GEN_880; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_882 = 8'h72 == io_in_3 ? 8'hcf : _GEN_881; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_883 = 8'h73 == io_in_3 ? 8'hc6 : _GEN_882; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_884 = 8'h74 == io_in_3 ? 8'hf9 : _GEN_883; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_885 = 8'h75 == io_in_3 ? 8'hf0 : _GEN_884; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_886 = 8'h76 == io_in_3 ? 8'heb : _GEN_885; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_887 = 8'h77 == io_in_3 ? 8'he2 : _GEN_886; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_888 = 8'h78 == io_in_3 ? 8'h95 : _GEN_887; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_889 = 8'h79 == io_in_3 ? 8'h9c : _GEN_888; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_890 = 8'h7a == io_in_3 ? 8'h87 : _GEN_889; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_891 = 8'h7b == io_in_3 ? 8'h8e : _GEN_890; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_892 = 8'h7c == io_in_3 ? 8'hb1 : _GEN_891; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_893 = 8'h7d == io_in_3 ? 8'hb8 : _GEN_892; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_894 = 8'h7e == io_in_3 ? 8'ha3 : _GEN_893; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_895 = 8'h7f == io_in_3 ? 8'haa : _GEN_894; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_896 = 8'h80 == io_in_3 ? 8'hec : _GEN_895; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_897 = 8'h81 == io_in_3 ? 8'he5 : _GEN_896; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_898 = 8'h82 == io_in_3 ? 8'hfe : _GEN_897; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_899 = 8'h83 == io_in_3 ? 8'hf7 : _GEN_898; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_900 = 8'h84 == io_in_3 ? 8'hc8 : _GEN_899; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_901 = 8'h85 == io_in_3 ? 8'hc1 : _GEN_900; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_902 = 8'h86 == io_in_3 ? 8'hda : _GEN_901; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_903 = 8'h87 == io_in_3 ? 8'hd3 : _GEN_902; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_904 = 8'h88 == io_in_3 ? 8'ha4 : _GEN_903; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_905 = 8'h89 == io_in_3 ? 8'had : _GEN_904; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_906 = 8'h8a == io_in_3 ? 8'hb6 : _GEN_905; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_907 = 8'h8b == io_in_3 ? 8'hbf : _GEN_906; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_908 = 8'h8c == io_in_3 ? 8'h80 : _GEN_907; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_909 = 8'h8d == io_in_3 ? 8'h89 : _GEN_908; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_910 = 8'h8e == io_in_3 ? 8'h92 : _GEN_909; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_911 = 8'h8f == io_in_3 ? 8'h9b : _GEN_910; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_912 = 8'h90 == io_in_3 ? 8'h7c : _GEN_911; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_913 = 8'h91 == io_in_3 ? 8'h75 : _GEN_912; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_914 = 8'h92 == io_in_3 ? 8'h6e : _GEN_913; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_915 = 8'h93 == io_in_3 ? 8'h67 : _GEN_914; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_916 = 8'h94 == io_in_3 ? 8'h58 : _GEN_915; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_917 = 8'h95 == io_in_3 ? 8'h51 : _GEN_916; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_918 = 8'h96 == io_in_3 ? 8'h4a : _GEN_917; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_919 = 8'h97 == io_in_3 ? 8'h43 : _GEN_918; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_920 = 8'h98 == io_in_3 ? 8'h34 : _GEN_919; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_921 = 8'h99 == io_in_3 ? 8'h3d : _GEN_920; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_922 = 8'h9a == io_in_3 ? 8'h26 : _GEN_921; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_923 = 8'h9b == io_in_3 ? 8'h2f : _GEN_922; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_924 = 8'h9c == io_in_3 ? 8'h10 : _GEN_923; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_925 = 8'h9d == io_in_3 ? 8'h19 : _GEN_924; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_926 = 8'h9e == io_in_3 ? 8'h2 : _GEN_925; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_927 = 8'h9f == io_in_3 ? 8'hb : _GEN_926; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_928 = 8'ha0 == io_in_3 ? 8'hd7 : _GEN_927; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_929 = 8'ha1 == io_in_3 ? 8'hde : _GEN_928; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_930 = 8'ha2 == io_in_3 ? 8'hc5 : _GEN_929; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_931 = 8'ha3 == io_in_3 ? 8'hcc : _GEN_930; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_932 = 8'ha4 == io_in_3 ? 8'hf3 : _GEN_931; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_933 = 8'ha5 == io_in_3 ? 8'hfa : _GEN_932; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_934 = 8'ha6 == io_in_3 ? 8'he1 : _GEN_933; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_935 = 8'ha7 == io_in_3 ? 8'he8 : _GEN_934; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_936 = 8'ha8 == io_in_3 ? 8'h9f : _GEN_935; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_937 = 8'ha9 == io_in_3 ? 8'h96 : _GEN_936; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_938 = 8'haa == io_in_3 ? 8'h8d : _GEN_937; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_939 = 8'hab == io_in_3 ? 8'h84 : _GEN_938; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_940 = 8'hac == io_in_3 ? 8'hbb : _GEN_939; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_941 = 8'had == io_in_3 ? 8'hb2 : _GEN_940; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_942 = 8'hae == io_in_3 ? 8'ha9 : _GEN_941; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_943 = 8'haf == io_in_3 ? 8'ha0 : _GEN_942; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_944 = 8'hb0 == io_in_3 ? 8'h47 : _GEN_943; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_945 = 8'hb1 == io_in_3 ? 8'h4e : _GEN_944; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_946 = 8'hb2 == io_in_3 ? 8'h55 : _GEN_945; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_947 = 8'hb3 == io_in_3 ? 8'h5c : _GEN_946; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_948 = 8'hb4 == io_in_3 ? 8'h63 : _GEN_947; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_949 = 8'hb5 == io_in_3 ? 8'h6a : _GEN_948; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_950 = 8'hb6 == io_in_3 ? 8'h71 : _GEN_949; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_951 = 8'hb7 == io_in_3 ? 8'h78 : _GEN_950; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_952 = 8'hb8 == io_in_3 ? 8'hf : _GEN_951; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_953 = 8'hb9 == io_in_3 ? 8'h6 : _GEN_952; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_954 = 8'hba == io_in_3 ? 8'h1d : _GEN_953; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_955 = 8'hbb == io_in_3 ? 8'h14 : _GEN_954; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_956 = 8'hbc == io_in_3 ? 8'h2b : _GEN_955; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_957 = 8'hbd == io_in_3 ? 8'h22 : _GEN_956; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_958 = 8'hbe == io_in_3 ? 8'h39 : _GEN_957; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_959 = 8'hbf == io_in_3 ? 8'h30 : _GEN_958; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_960 = 8'hc0 == io_in_3 ? 8'h9a : _GEN_959; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_961 = 8'hc1 == io_in_3 ? 8'h93 : _GEN_960; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_962 = 8'hc2 == io_in_3 ? 8'h88 : _GEN_961; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_963 = 8'hc3 == io_in_3 ? 8'h81 : _GEN_962; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_964 = 8'hc4 == io_in_3 ? 8'hbe : _GEN_963; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_965 = 8'hc5 == io_in_3 ? 8'hb7 : _GEN_964; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_966 = 8'hc6 == io_in_3 ? 8'hac : _GEN_965; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_967 = 8'hc7 == io_in_3 ? 8'ha5 : _GEN_966; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_968 = 8'hc8 == io_in_3 ? 8'hd2 : _GEN_967; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_969 = 8'hc9 == io_in_3 ? 8'hdb : _GEN_968; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_970 = 8'hca == io_in_3 ? 8'hc0 : _GEN_969; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_971 = 8'hcb == io_in_3 ? 8'hc9 : _GEN_970; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_972 = 8'hcc == io_in_3 ? 8'hf6 : _GEN_971; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_973 = 8'hcd == io_in_3 ? 8'hff : _GEN_972; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_974 = 8'hce == io_in_3 ? 8'he4 : _GEN_973; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_975 = 8'hcf == io_in_3 ? 8'hed : _GEN_974; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_976 = 8'hd0 == io_in_3 ? 8'ha : _GEN_975; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_977 = 8'hd1 == io_in_3 ? 8'h3 : _GEN_976; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_978 = 8'hd2 == io_in_3 ? 8'h18 : _GEN_977; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_979 = 8'hd3 == io_in_3 ? 8'h11 : _GEN_978; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_980 = 8'hd4 == io_in_3 ? 8'h2e : _GEN_979; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_981 = 8'hd5 == io_in_3 ? 8'h27 : _GEN_980; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_982 = 8'hd6 == io_in_3 ? 8'h3c : _GEN_981; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_983 = 8'hd7 == io_in_3 ? 8'h35 : _GEN_982; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_984 = 8'hd8 == io_in_3 ? 8'h42 : _GEN_983; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_985 = 8'hd9 == io_in_3 ? 8'h4b : _GEN_984; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_986 = 8'hda == io_in_3 ? 8'h50 : _GEN_985; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_987 = 8'hdb == io_in_3 ? 8'h59 : _GEN_986; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_988 = 8'hdc == io_in_3 ? 8'h66 : _GEN_987; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_989 = 8'hdd == io_in_3 ? 8'h6f : _GEN_988; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_990 = 8'hde == io_in_3 ? 8'h74 : _GEN_989; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_991 = 8'hdf == io_in_3 ? 8'h7d : _GEN_990; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_992 = 8'he0 == io_in_3 ? 8'ha1 : _GEN_991; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_993 = 8'he1 == io_in_3 ? 8'ha8 : _GEN_992; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_994 = 8'he2 == io_in_3 ? 8'hb3 : _GEN_993; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_995 = 8'he3 == io_in_3 ? 8'hba : _GEN_994; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_996 = 8'he4 == io_in_3 ? 8'h85 : _GEN_995; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_997 = 8'he5 == io_in_3 ? 8'h8c : _GEN_996; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_998 = 8'he6 == io_in_3 ? 8'h97 : _GEN_997; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_999 = 8'he7 == io_in_3 ? 8'h9e : _GEN_998; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1000 = 8'he8 == io_in_3 ? 8'he9 : _GEN_999; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1001 = 8'he9 == io_in_3 ? 8'he0 : _GEN_1000; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1002 = 8'hea == io_in_3 ? 8'hfb : _GEN_1001; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1003 = 8'heb == io_in_3 ? 8'hf2 : _GEN_1002; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1004 = 8'hec == io_in_3 ? 8'hcd : _GEN_1003; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1005 = 8'hed == io_in_3 ? 8'hc4 : _GEN_1004; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1006 = 8'hee == io_in_3 ? 8'hdf : _GEN_1005; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1007 = 8'hef == io_in_3 ? 8'hd6 : _GEN_1006; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1008 = 8'hf0 == io_in_3 ? 8'h31 : _GEN_1007; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1009 = 8'hf1 == io_in_3 ? 8'h38 : _GEN_1008; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1010 = 8'hf2 == io_in_3 ? 8'h23 : _GEN_1009; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1011 = 8'hf3 == io_in_3 ? 8'h2a : _GEN_1010; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1012 = 8'hf4 == io_in_3 ? 8'h15 : _GEN_1011; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1013 = 8'hf5 == io_in_3 ? 8'h1c : _GEN_1012; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1014 = 8'hf6 == io_in_3 ? 8'h7 : _GEN_1013; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1015 = 8'hf7 == io_in_3 ? 8'he : _GEN_1014; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1016 = 8'hf8 == io_in_3 ? 8'h79 : _GEN_1015; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1017 = 8'hf9 == io_in_3 ? 8'h70 : _GEN_1016; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1018 = 8'hfa == io_in_3 ? 8'h6b : _GEN_1017; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1019 = 8'hfb == io_in_3 ? 8'h62 : _GEN_1018; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1020 = 8'hfc == io_in_3 ? 8'h5d : _GEN_1019; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1021 = 8'hfd == io_in_3 ? 8'h54 : _GEN_1020; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1022 = 8'hfe == io_in_3 ? 8'h4f : _GEN_1021; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1023 = 8'hff == io_in_3 ? 8'h46 : _GEN_1022; // @[AES_PipelinedElasticBuffer.scala 591:68 AES_PipelinedElasticBuffer.scala 591:68]
  wire [7:0] _GEN_1025 = 8'h1 == io_in_0 ? 8'h9 : 8'h0; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1026 = 8'h2 == io_in_0 ? 8'h12 : _GEN_1025; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1027 = 8'h3 == io_in_0 ? 8'h1b : _GEN_1026; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1028 = 8'h4 == io_in_0 ? 8'h24 : _GEN_1027; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1029 = 8'h5 == io_in_0 ? 8'h2d : _GEN_1028; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1030 = 8'h6 == io_in_0 ? 8'h36 : _GEN_1029; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1031 = 8'h7 == io_in_0 ? 8'h3f : _GEN_1030; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1032 = 8'h8 == io_in_0 ? 8'h48 : _GEN_1031; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1033 = 8'h9 == io_in_0 ? 8'h41 : _GEN_1032; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1034 = 8'ha == io_in_0 ? 8'h5a : _GEN_1033; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1035 = 8'hb == io_in_0 ? 8'h53 : _GEN_1034; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1036 = 8'hc == io_in_0 ? 8'h6c : _GEN_1035; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1037 = 8'hd == io_in_0 ? 8'h65 : _GEN_1036; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1038 = 8'he == io_in_0 ? 8'h7e : _GEN_1037; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1039 = 8'hf == io_in_0 ? 8'h77 : _GEN_1038; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1040 = 8'h10 == io_in_0 ? 8'h90 : _GEN_1039; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1041 = 8'h11 == io_in_0 ? 8'h99 : _GEN_1040; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1042 = 8'h12 == io_in_0 ? 8'h82 : _GEN_1041; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1043 = 8'h13 == io_in_0 ? 8'h8b : _GEN_1042; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1044 = 8'h14 == io_in_0 ? 8'hb4 : _GEN_1043; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1045 = 8'h15 == io_in_0 ? 8'hbd : _GEN_1044; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1046 = 8'h16 == io_in_0 ? 8'ha6 : _GEN_1045; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1047 = 8'h17 == io_in_0 ? 8'haf : _GEN_1046; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1048 = 8'h18 == io_in_0 ? 8'hd8 : _GEN_1047; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1049 = 8'h19 == io_in_0 ? 8'hd1 : _GEN_1048; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1050 = 8'h1a == io_in_0 ? 8'hca : _GEN_1049; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1051 = 8'h1b == io_in_0 ? 8'hc3 : _GEN_1050; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1052 = 8'h1c == io_in_0 ? 8'hfc : _GEN_1051; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1053 = 8'h1d == io_in_0 ? 8'hf5 : _GEN_1052; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1054 = 8'h1e == io_in_0 ? 8'hee : _GEN_1053; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1055 = 8'h1f == io_in_0 ? 8'he7 : _GEN_1054; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1056 = 8'h20 == io_in_0 ? 8'h3b : _GEN_1055; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1057 = 8'h21 == io_in_0 ? 8'h32 : _GEN_1056; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1058 = 8'h22 == io_in_0 ? 8'h29 : _GEN_1057; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1059 = 8'h23 == io_in_0 ? 8'h20 : _GEN_1058; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1060 = 8'h24 == io_in_0 ? 8'h1f : _GEN_1059; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1061 = 8'h25 == io_in_0 ? 8'h16 : _GEN_1060; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1062 = 8'h26 == io_in_0 ? 8'hd : _GEN_1061; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1063 = 8'h27 == io_in_0 ? 8'h4 : _GEN_1062; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1064 = 8'h28 == io_in_0 ? 8'h73 : _GEN_1063; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1065 = 8'h29 == io_in_0 ? 8'h7a : _GEN_1064; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1066 = 8'h2a == io_in_0 ? 8'h61 : _GEN_1065; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1067 = 8'h2b == io_in_0 ? 8'h68 : _GEN_1066; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1068 = 8'h2c == io_in_0 ? 8'h57 : _GEN_1067; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1069 = 8'h2d == io_in_0 ? 8'h5e : _GEN_1068; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1070 = 8'h2e == io_in_0 ? 8'h45 : _GEN_1069; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1071 = 8'h2f == io_in_0 ? 8'h4c : _GEN_1070; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1072 = 8'h30 == io_in_0 ? 8'hab : _GEN_1071; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1073 = 8'h31 == io_in_0 ? 8'ha2 : _GEN_1072; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1074 = 8'h32 == io_in_0 ? 8'hb9 : _GEN_1073; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1075 = 8'h33 == io_in_0 ? 8'hb0 : _GEN_1074; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1076 = 8'h34 == io_in_0 ? 8'h8f : _GEN_1075; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1077 = 8'h35 == io_in_0 ? 8'h86 : _GEN_1076; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1078 = 8'h36 == io_in_0 ? 8'h9d : _GEN_1077; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1079 = 8'h37 == io_in_0 ? 8'h94 : _GEN_1078; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1080 = 8'h38 == io_in_0 ? 8'he3 : _GEN_1079; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1081 = 8'h39 == io_in_0 ? 8'hea : _GEN_1080; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1082 = 8'h3a == io_in_0 ? 8'hf1 : _GEN_1081; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1083 = 8'h3b == io_in_0 ? 8'hf8 : _GEN_1082; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1084 = 8'h3c == io_in_0 ? 8'hc7 : _GEN_1083; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1085 = 8'h3d == io_in_0 ? 8'hce : _GEN_1084; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1086 = 8'h3e == io_in_0 ? 8'hd5 : _GEN_1085; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1087 = 8'h3f == io_in_0 ? 8'hdc : _GEN_1086; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1088 = 8'h40 == io_in_0 ? 8'h76 : _GEN_1087; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1089 = 8'h41 == io_in_0 ? 8'h7f : _GEN_1088; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1090 = 8'h42 == io_in_0 ? 8'h64 : _GEN_1089; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1091 = 8'h43 == io_in_0 ? 8'h6d : _GEN_1090; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1092 = 8'h44 == io_in_0 ? 8'h52 : _GEN_1091; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1093 = 8'h45 == io_in_0 ? 8'h5b : _GEN_1092; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1094 = 8'h46 == io_in_0 ? 8'h40 : _GEN_1093; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1095 = 8'h47 == io_in_0 ? 8'h49 : _GEN_1094; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1096 = 8'h48 == io_in_0 ? 8'h3e : _GEN_1095; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1097 = 8'h49 == io_in_0 ? 8'h37 : _GEN_1096; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1098 = 8'h4a == io_in_0 ? 8'h2c : _GEN_1097; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1099 = 8'h4b == io_in_0 ? 8'h25 : _GEN_1098; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1100 = 8'h4c == io_in_0 ? 8'h1a : _GEN_1099; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1101 = 8'h4d == io_in_0 ? 8'h13 : _GEN_1100; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1102 = 8'h4e == io_in_0 ? 8'h8 : _GEN_1101; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1103 = 8'h4f == io_in_0 ? 8'h1 : _GEN_1102; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1104 = 8'h50 == io_in_0 ? 8'he6 : _GEN_1103; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1105 = 8'h51 == io_in_0 ? 8'hef : _GEN_1104; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1106 = 8'h52 == io_in_0 ? 8'hf4 : _GEN_1105; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1107 = 8'h53 == io_in_0 ? 8'hfd : _GEN_1106; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1108 = 8'h54 == io_in_0 ? 8'hc2 : _GEN_1107; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1109 = 8'h55 == io_in_0 ? 8'hcb : _GEN_1108; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1110 = 8'h56 == io_in_0 ? 8'hd0 : _GEN_1109; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1111 = 8'h57 == io_in_0 ? 8'hd9 : _GEN_1110; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1112 = 8'h58 == io_in_0 ? 8'hae : _GEN_1111; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1113 = 8'h59 == io_in_0 ? 8'ha7 : _GEN_1112; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1114 = 8'h5a == io_in_0 ? 8'hbc : _GEN_1113; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1115 = 8'h5b == io_in_0 ? 8'hb5 : _GEN_1114; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1116 = 8'h5c == io_in_0 ? 8'h8a : _GEN_1115; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1117 = 8'h5d == io_in_0 ? 8'h83 : _GEN_1116; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1118 = 8'h5e == io_in_0 ? 8'h98 : _GEN_1117; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1119 = 8'h5f == io_in_0 ? 8'h91 : _GEN_1118; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1120 = 8'h60 == io_in_0 ? 8'h4d : _GEN_1119; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1121 = 8'h61 == io_in_0 ? 8'h44 : _GEN_1120; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1122 = 8'h62 == io_in_0 ? 8'h5f : _GEN_1121; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1123 = 8'h63 == io_in_0 ? 8'h56 : _GEN_1122; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1124 = 8'h64 == io_in_0 ? 8'h69 : _GEN_1123; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1125 = 8'h65 == io_in_0 ? 8'h60 : _GEN_1124; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1126 = 8'h66 == io_in_0 ? 8'h7b : _GEN_1125; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1127 = 8'h67 == io_in_0 ? 8'h72 : _GEN_1126; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1128 = 8'h68 == io_in_0 ? 8'h5 : _GEN_1127; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1129 = 8'h69 == io_in_0 ? 8'hc : _GEN_1128; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1130 = 8'h6a == io_in_0 ? 8'h17 : _GEN_1129; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1131 = 8'h6b == io_in_0 ? 8'h1e : _GEN_1130; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1132 = 8'h6c == io_in_0 ? 8'h21 : _GEN_1131; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1133 = 8'h6d == io_in_0 ? 8'h28 : _GEN_1132; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1134 = 8'h6e == io_in_0 ? 8'h33 : _GEN_1133; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1135 = 8'h6f == io_in_0 ? 8'h3a : _GEN_1134; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1136 = 8'h70 == io_in_0 ? 8'hdd : _GEN_1135; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1137 = 8'h71 == io_in_0 ? 8'hd4 : _GEN_1136; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1138 = 8'h72 == io_in_0 ? 8'hcf : _GEN_1137; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1139 = 8'h73 == io_in_0 ? 8'hc6 : _GEN_1138; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1140 = 8'h74 == io_in_0 ? 8'hf9 : _GEN_1139; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1141 = 8'h75 == io_in_0 ? 8'hf0 : _GEN_1140; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1142 = 8'h76 == io_in_0 ? 8'heb : _GEN_1141; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1143 = 8'h77 == io_in_0 ? 8'he2 : _GEN_1142; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1144 = 8'h78 == io_in_0 ? 8'h95 : _GEN_1143; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1145 = 8'h79 == io_in_0 ? 8'h9c : _GEN_1144; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1146 = 8'h7a == io_in_0 ? 8'h87 : _GEN_1145; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1147 = 8'h7b == io_in_0 ? 8'h8e : _GEN_1146; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1148 = 8'h7c == io_in_0 ? 8'hb1 : _GEN_1147; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1149 = 8'h7d == io_in_0 ? 8'hb8 : _GEN_1148; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1150 = 8'h7e == io_in_0 ? 8'ha3 : _GEN_1149; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1151 = 8'h7f == io_in_0 ? 8'haa : _GEN_1150; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1152 = 8'h80 == io_in_0 ? 8'hec : _GEN_1151; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1153 = 8'h81 == io_in_0 ? 8'he5 : _GEN_1152; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1154 = 8'h82 == io_in_0 ? 8'hfe : _GEN_1153; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1155 = 8'h83 == io_in_0 ? 8'hf7 : _GEN_1154; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1156 = 8'h84 == io_in_0 ? 8'hc8 : _GEN_1155; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1157 = 8'h85 == io_in_0 ? 8'hc1 : _GEN_1156; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1158 = 8'h86 == io_in_0 ? 8'hda : _GEN_1157; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1159 = 8'h87 == io_in_0 ? 8'hd3 : _GEN_1158; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1160 = 8'h88 == io_in_0 ? 8'ha4 : _GEN_1159; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1161 = 8'h89 == io_in_0 ? 8'had : _GEN_1160; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1162 = 8'h8a == io_in_0 ? 8'hb6 : _GEN_1161; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1163 = 8'h8b == io_in_0 ? 8'hbf : _GEN_1162; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1164 = 8'h8c == io_in_0 ? 8'h80 : _GEN_1163; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1165 = 8'h8d == io_in_0 ? 8'h89 : _GEN_1164; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1166 = 8'h8e == io_in_0 ? 8'h92 : _GEN_1165; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1167 = 8'h8f == io_in_0 ? 8'h9b : _GEN_1166; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1168 = 8'h90 == io_in_0 ? 8'h7c : _GEN_1167; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1169 = 8'h91 == io_in_0 ? 8'h75 : _GEN_1168; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1170 = 8'h92 == io_in_0 ? 8'h6e : _GEN_1169; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1171 = 8'h93 == io_in_0 ? 8'h67 : _GEN_1170; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1172 = 8'h94 == io_in_0 ? 8'h58 : _GEN_1171; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1173 = 8'h95 == io_in_0 ? 8'h51 : _GEN_1172; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1174 = 8'h96 == io_in_0 ? 8'h4a : _GEN_1173; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1175 = 8'h97 == io_in_0 ? 8'h43 : _GEN_1174; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1176 = 8'h98 == io_in_0 ? 8'h34 : _GEN_1175; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1177 = 8'h99 == io_in_0 ? 8'h3d : _GEN_1176; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1178 = 8'h9a == io_in_0 ? 8'h26 : _GEN_1177; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1179 = 8'h9b == io_in_0 ? 8'h2f : _GEN_1178; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1180 = 8'h9c == io_in_0 ? 8'h10 : _GEN_1179; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1181 = 8'h9d == io_in_0 ? 8'h19 : _GEN_1180; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1182 = 8'h9e == io_in_0 ? 8'h2 : _GEN_1181; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1183 = 8'h9f == io_in_0 ? 8'hb : _GEN_1182; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1184 = 8'ha0 == io_in_0 ? 8'hd7 : _GEN_1183; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1185 = 8'ha1 == io_in_0 ? 8'hde : _GEN_1184; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1186 = 8'ha2 == io_in_0 ? 8'hc5 : _GEN_1185; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1187 = 8'ha3 == io_in_0 ? 8'hcc : _GEN_1186; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1188 = 8'ha4 == io_in_0 ? 8'hf3 : _GEN_1187; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1189 = 8'ha5 == io_in_0 ? 8'hfa : _GEN_1188; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1190 = 8'ha6 == io_in_0 ? 8'he1 : _GEN_1189; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1191 = 8'ha7 == io_in_0 ? 8'he8 : _GEN_1190; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1192 = 8'ha8 == io_in_0 ? 8'h9f : _GEN_1191; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1193 = 8'ha9 == io_in_0 ? 8'h96 : _GEN_1192; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1194 = 8'haa == io_in_0 ? 8'h8d : _GEN_1193; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1195 = 8'hab == io_in_0 ? 8'h84 : _GEN_1194; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1196 = 8'hac == io_in_0 ? 8'hbb : _GEN_1195; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1197 = 8'had == io_in_0 ? 8'hb2 : _GEN_1196; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1198 = 8'hae == io_in_0 ? 8'ha9 : _GEN_1197; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1199 = 8'haf == io_in_0 ? 8'ha0 : _GEN_1198; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1200 = 8'hb0 == io_in_0 ? 8'h47 : _GEN_1199; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1201 = 8'hb1 == io_in_0 ? 8'h4e : _GEN_1200; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1202 = 8'hb2 == io_in_0 ? 8'h55 : _GEN_1201; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1203 = 8'hb3 == io_in_0 ? 8'h5c : _GEN_1202; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1204 = 8'hb4 == io_in_0 ? 8'h63 : _GEN_1203; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1205 = 8'hb5 == io_in_0 ? 8'h6a : _GEN_1204; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1206 = 8'hb6 == io_in_0 ? 8'h71 : _GEN_1205; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1207 = 8'hb7 == io_in_0 ? 8'h78 : _GEN_1206; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1208 = 8'hb8 == io_in_0 ? 8'hf : _GEN_1207; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1209 = 8'hb9 == io_in_0 ? 8'h6 : _GEN_1208; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1210 = 8'hba == io_in_0 ? 8'h1d : _GEN_1209; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1211 = 8'hbb == io_in_0 ? 8'h14 : _GEN_1210; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1212 = 8'hbc == io_in_0 ? 8'h2b : _GEN_1211; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1213 = 8'hbd == io_in_0 ? 8'h22 : _GEN_1212; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1214 = 8'hbe == io_in_0 ? 8'h39 : _GEN_1213; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1215 = 8'hbf == io_in_0 ? 8'h30 : _GEN_1214; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1216 = 8'hc0 == io_in_0 ? 8'h9a : _GEN_1215; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1217 = 8'hc1 == io_in_0 ? 8'h93 : _GEN_1216; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1218 = 8'hc2 == io_in_0 ? 8'h88 : _GEN_1217; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1219 = 8'hc3 == io_in_0 ? 8'h81 : _GEN_1218; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1220 = 8'hc4 == io_in_0 ? 8'hbe : _GEN_1219; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1221 = 8'hc5 == io_in_0 ? 8'hb7 : _GEN_1220; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1222 = 8'hc6 == io_in_0 ? 8'hac : _GEN_1221; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1223 = 8'hc7 == io_in_0 ? 8'ha5 : _GEN_1222; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1224 = 8'hc8 == io_in_0 ? 8'hd2 : _GEN_1223; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1225 = 8'hc9 == io_in_0 ? 8'hdb : _GEN_1224; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1226 = 8'hca == io_in_0 ? 8'hc0 : _GEN_1225; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1227 = 8'hcb == io_in_0 ? 8'hc9 : _GEN_1226; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1228 = 8'hcc == io_in_0 ? 8'hf6 : _GEN_1227; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1229 = 8'hcd == io_in_0 ? 8'hff : _GEN_1228; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1230 = 8'hce == io_in_0 ? 8'he4 : _GEN_1229; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1231 = 8'hcf == io_in_0 ? 8'hed : _GEN_1230; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1232 = 8'hd0 == io_in_0 ? 8'ha : _GEN_1231; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1233 = 8'hd1 == io_in_0 ? 8'h3 : _GEN_1232; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1234 = 8'hd2 == io_in_0 ? 8'h18 : _GEN_1233; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1235 = 8'hd3 == io_in_0 ? 8'h11 : _GEN_1234; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1236 = 8'hd4 == io_in_0 ? 8'h2e : _GEN_1235; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1237 = 8'hd5 == io_in_0 ? 8'h27 : _GEN_1236; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1238 = 8'hd6 == io_in_0 ? 8'h3c : _GEN_1237; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1239 = 8'hd7 == io_in_0 ? 8'h35 : _GEN_1238; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1240 = 8'hd8 == io_in_0 ? 8'h42 : _GEN_1239; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1241 = 8'hd9 == io_in_0 ? 8'h4b : _GEN_1240; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1242 = 8'hda == io_in_0 ? 8'h50 : _GEN_1241; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1243 = 8'hdb == io_in_0 ? 8'h59 : _GEN_1242; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1244 = 8'hdc == io_in_0 ? 8'h66 : _GEN_1243; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1245 = 8'hdd == io_in_0 ? 8'h6f : _GEN_1244; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1246 = 8'hde == io_in_0 ? 8'h74 : _GEN_1245; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1247 = 8'hdf == io_in_0 ? 8'h7d : _GEN_1246; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1248 = 8'he0 == io_in_0 ? 8'ha1 : _GEN_1247; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1249 = 8'he1 == io_in_0 ? 8'ha8 : _GEN_1248; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1250 = 8'he2 == io_in_0 ? 8'hb3 : _GEN_1249; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1251 = 8'he3 == io_in_0 ? 8'hba : _GEN_1250; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1252 = 8'he4 == io_in_0 ? 8'h85 : _GEN_1251; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1253 = 8'he5 == io_in_0 ? 8'h8c : _GEN_1252; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1254 = 8'he6 == io_in_0 ? 8'h97 : _GEN_1253; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1255 = 8'he7 == io_in_0 ? 8'h9e : _GEN_1254; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1256 = 8'he8 == io_in_0 ? 8'he9 : _GEN_1255; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1257 = 8'he9 == io_in_0 ? 8'he0 : _GEN_1256; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1258 = 8'hea == io_in_0 ? 8'hfb : _GEN_1257; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1259 = 8'heb == io_in_0 ? 8'hf2 : _GEN_1258; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1260 = 8'hec == io_in_0 ? 8'hcd : _GEN_1259; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1261 = 8'hed == io_in_0 ? 8'hc4 : _GEN_1260; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1262 = 8'hee == io_in_0 ? 8'hdf : _GEN_1261; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1263 = 8'hef == io_in_0 ? 8'hd6 : _GEN_1262; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1264 = 8'hf0 == io_in_0 ? 8'h31 : _GEN_1263; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1265 = 8'hf1 == io_in_0 ? 8'h38 : _GEN_1264; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1266 = 8'hf2 == io_in_0 ? 8'h23 : _GEN_1265; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1267 = 8'hf3 == io_in_0 ? 8'h2a : _GEN_1266; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1268 = 8'hf4 == io_in_0 ? 8'h15 : _GEN_1267; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1269 = 8'hf5 == io_in_0 ? 8'h1c : _GEN_1268; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1270 = 8'hf6 == io_in_0 ? 8'h7 : _GEN_1269; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1271 = 8'hf7 == io_in_0 ? 8'he : _GEN_1270; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1272 = 8'hf8 == io_in_0 ? 8'h79 : _GEN_1271; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1273 = 8'hf9 == io_in_0 ? 8'h70 : _GEN_1272; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1274 = 8'hfa == io_in_0 ? 8'h6b : _GEN_1273; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1275 = 8'hfb == io_in_0 ? 8'h62 : _GEN_1274; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1276 = 8'hfc == io_in_0 ? 8'h5d : _GEN_1275; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1277 = 8'hfd == io_in_0 ? 8'h54 : _GEN_1276; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1278 = 8'hfe == io_in_0 ? 8'h4f : _GEN_1277; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1279 = 8'hff == io_in_0 ? 8'h46 : _GEN_1278; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1281 = 8'h1 == io_in_1 ? 8'he : 8'h0; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1282 = 8'h2 == io_in_1 ? 8'h1c : _GEN_1281; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1283 = 8'h3 == io_in_1 ? 8'h12 : _GEN_1282; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1284 = 8'h4 == io_in_1 ? 8'h38 : _GEN_1283; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1285 = 8'h5 == io_in_1 ? 8'h36 : _GEN_1284; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1286 = 8'h6 == io_in_1 ? 8'h24 : _GEN_1285; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1287 = 8'h7 == io_in_1 ? 8'h2a : _GEN_1286; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1288 = 8'h8 == io_in_1 ? 8'h70 : _GEN_1287; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1289 = 8'h9 == io_in_1 ? 8'h7e : _GEN_1288; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1290 = 8'ha == io_in_1 ? 8'h6c : _GEN_1289; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1291 = 8'hb == io_in_1 ? 8'h62 : _GEN_1290; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1292 = 8'hc == io_in_1 ? 8'h48 : _GEN_1291; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1293 = 8'hd == io_in_1 ? 8'h46 : _GEN_1292; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1294 = 8'he == io_in_1 ? 8'h54 : _GEN_1293; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1295 = 8'hf == io_in_1 ? 8'h5a : _GEN_1294; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1296 = 8'h10 == io_in_1 ? 8'he0 : _GEN_1295; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1297 = 8'h11 == io_in_1 ? 8'hee : _GEN_1296; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1298 = 8'h12 == io_in_1 ? 8'hfc : _GEN_1297; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1299 = 8'h13 == io_in_1 ? 8'hf2 : _GEN_1298; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1300 = 8'h14 == io_in_1 ? 8'hd8 : _GEN_1299; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1301 = 8'h15 == io_in_1 ? 8'hd6 : _GEN_1300; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1302 = 8'h16 == io_in_1 ? 8'hc4 : _GEN_1301; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1303 = 8'h17 == io_in_1 ? 8'hca : _GEN_1302; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1304 = 8'h18 == io_in_1 ? 8'h90 : _GEN_1303; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1305 = 8'h19 == io_in_1 ? 8'h9e : _GEN_1304; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1306 = 8'h1a == io_in_1 ? 8'h8c : _GEN_1305; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1307 = 8'h1b == io_in_1 ? 8'h82 : _GEN_1306; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1308 = 8'h1c == io_in_1 ? 8'ha8 : _GEN_1307; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1309 = 8'h1d == io_in_1 ? 8'ha6 : _GEN_1308; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1310 = 8'h1e == io_in_1 ? 8'hb4 : _GEN_1309; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1311 = 8'h1f == io_in_1 ? 8'hba : _GEN_1310; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1312 = 8'h20 == io_in_1 ? 8'hdb : _GEN_1311; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1313 = 8'h21 == io_in_1 ? 8'hd5 : _GEN_1312; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1314 = 8'h22 == io_in_1 ? 8'hc7 : _GEN_1313; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1315 = 8'h23 == io_in_1 ? 8'hc9 : _GEN_1314; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1316 = 8'h24 == io_in_1 ? 8'he3 : _GEN_1315; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1317 = 8'h25 == io_in_1 ? 8'hed : _GEN_1316; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1318 = 8'h26 == io_in_1 ? 8'hff : _GEN_1317; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1319 = 8'h27 == io_in_1 ? 8'hf1 : _GEN_1318; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1320 = 8'h28 == io_in_1 ? 8'hab : _GEN_1319; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1321 = 8'h29 == io_in_1 ? 8'ha5 : _GEN_1320; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1322 = 8'h2a == io_in_1 ? 8'hb7 : _GEN_1321; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1323 = 8'h2b == io_in_1 ? 8'hb9 : _GEN_1322; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1324 = 8'h2c == io_in_1 ? 8'h93 : _GEN_1323; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1325 = 8'h2d == io_in_1 ? 8'h9d : _GEN_1324; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1326 = 8'h2e == io_in_1 ? 8'h8f : _GEN_1325; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1327 = 8'h2f == io_in_1 ? 8'h81 : _GEN_1326; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1328 = 8'h30 == io_in_1 ? 8'h3b : _GEN_1327; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1329 = 8'h31 == io_in_1 ? 8'h35 : _GEN_1328; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1330 = 8'h32 == io_in_1 ? 8'h27 : _GEN_1329; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1331 = 8'h33 == io_in_1 ? 8'h29 : _GEN_1330; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1332 = 8'h34 == io_in_1 ? 8'h3 : _GEN_1331; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1333 = 8'h35 == io_in_1 ? 8'hd : _GEN_1332; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1334 = 8'h36 == io_in_1 ? 8'h1f : _GEN_1333; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1335 = 8'h37 == io_in_1 ? 8'h11 : _GEN_1334; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1336 = 8'h38 == io_in_1 ? 8'h4b : _GEN_1335; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1337 = 8'h39 == io_in_1 ? 8'h45 : _GEN_1336; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1338 = 8'h3a == io_in_1 ? 8'h57 : _GEN_1337; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1339 = 8'h3b == io_in_1 ? 8'h59 : _GEN_1338; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1340 = 8'h3c == io_in_1 ? 8'h73 : _GEN_1339; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1341 = 8'h3d == io_in_1 ? 8'h7d : _GEN_1340; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1342 = 8'h3e == io_in_1 ? 8'h6f : _GEN_1341; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1343 = 8'h3f == io_in_1 ? 8'h61 : _GEN_1342; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1344 = 8'h40 == io_in_1 ? 8'had : _GEN_1343; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1345 = 8'h41 == io_in_1 ? 8'ha3 : _GEN_1344; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1346 = 8'h42 == io_in_1 ? 8'hb1 : _GEN_1345; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1347 = 8'h43 == io_in_1 ? 8'hbf : _GEN_1346; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1348 = 8'h44 == io_in_1 ? 8'h95 : _GEN_1347; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1349 = 8'h45 == io_in_1 ? 8'h9b : _GEN_1348; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1350 = 8'h46 == io_in_1 ? 8'h89 : _GEN_1349; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1351 = 8'h47 == io_in_1 ? 8'h87 : _GEN_1350; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1352 = 8'h48 == io_in_1 ? 8'hdd : _GEN_1351; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1353 = 8'h49 == io_in_1 ? 8'hd3 : _GEN_1352; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1354 = 8'h4a == io_in_1 ? 8'hc1 : _GEN_1353; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1355 = 8'h4b == io_in_1 ? 8'hcf : _GEN_1354; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1356 = 8'h4c == io_in_1 ? 8'he5 : _GEN_1355; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1357 = 8'h4d == io_in_1 ? 8'heb : _GEN_1356; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1358 = 8'h4e == io_in_1 ? 8'hf9 : _GEN_1357; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1359 = 8'h4f == io_in_1 ? 8'hf7 : _GEN_1358; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1360 = 8'h50 == io_in_1 ? 8'h4d : _GEN_1359; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1361 = 8'h51 == io_in_1 ? 8'h43 : _GEN_1360; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1362 = 8'h52 == io_in_1 ? 8'h51 : _GEN_1361; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1363 = 8'h53 == io_in_1 ? 8'h5f : _GEN_1362; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1364 = 8'h54 == io_in_1 ? 8'h75 : _GEN_1363; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1365 = 8'h55 == io_in_1 ? 8'h7b : _GEN_1364; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1366 = 8'h56 == io_in_1 ? 8'h69 : _GEN_1365; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1367 = 8'h57 == io_in_1 ? 8'h67 : _GEN_1366; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1368 = 8'h58 == io_in_1 ? 8'h3d : _GEN_1367; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1369 = 8'h59 == io_in_1 ? 8'h33 : _GEN_1368; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1370 = 8'h5a == io_in_1 ? 8'h21 : _GEN_1369; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1371 = 8'h5b == io_in_1 ? 8'h2f : _GEN_1370; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1372 = 8'h5c == io_in_1 ? 8'h5 : _GEN_1371; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1373 = 8'h5d == io_in_1 ? 8'hb : _GEN_1372; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1374 = 8'h5e == io_in_1 ? 8'h19 : _GEN_1373; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1375 = 8'h5f == io_in_1 ? 8'h17 : _GEN_1374; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1376 = 8'h60 == io_in_1 ? 8'h76 : _GEN_1375; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1377 = 8'h61 == io_in_1 ? 8'h78 : _GEN_1376; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1378 = 8'h62 == io_in_1 ? 8'h6a : _GEN_1377; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1379 = 8'h63 == io_in_1 ? 8'h64 : _GEN_1378; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1380 = 8'h64 == io_in_1 ? 8'h4e : _GEN_1379; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1381 = 8'h65 == io_in_1 ? 8'h40 : _GEN_1380; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1382 = 8'h66 == io_in_1 ? 8'h52 : _GEN_1381; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1383 = 8'h67 == io_in_1 ? 8'h5c : _GEN_1382; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1384 = 8'h68 == io_in_1 ? 8'h6 : _GEN_1383; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1385 = 8'h69 == io_in_1 ? 8'h8 : _GEN_1384; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1386 = 8'h6a == io_in_1 ? 8'h1a : _GEN_1385; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1387 = 8'h6b == io_in_1 ? 8'h14 : _GEN_1386; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1388 = 8'h6c == io_in_1 ? 8'h3e : _GEN_1387; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1389 = 8'h6d == io_in_1 ? 8'h30 : _GEN_1388; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1390 = 8'h6e == io_in_1 ? 8'h22 : _GEN_1389; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1391 = 8'h6f == io_in_1 ? 8'h2c : _GEN_1390; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1392 = 8'h70 == io_in_1 ? 8'h96 : _GEN_1391; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1393 = 8'h71 == io_in_1 ? 8'h98 : _GEN_1392; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1394 = 8'h72 == io_in_1 ? 8'h8a : _GEN_1393; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1395 = 8'h73 == io_in_1 ? 8'h84 : _GEN_1394; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1396 = 8'h74 == io_in_1 ? 8'hae : _GEN_1395; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1397 = 8'h75 == io_in_1 ? 8'ha0 : _GEN_1396; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1398 = 8'h76 == io_in_1 ? 8'hb2 : _GEN_1397; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1399 = 8'h77 == io_in_1 ? 8'hbc : _GEN_1398; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1400 = 8'h78 == io_in_1 ? 8'he6 : _GEN_1399; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1401 = 8'h79 == io_in_1 ? 8'he8 : _GEN_1400; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1402 = 8'h7a == io_in_1 ? 8'hfa : _GEN_1401; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1403 = 8'h7b == io_in_1 ? 8'hf4 : _GEN_1402; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1404 = 8'h7c == io_in_1 ? 8'hde : _GEN_1403; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1405 = 8'h7d == io_in_1 ? 8'hd0 : _GEN_1404; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1406 = 8'h7e == io_in_1 ? 8'hc2 : _GEN_1405; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1407 = 8'h7f == io_in_1 ? 8'hcc : _GEN_1406; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1408 = 8'h80 == io_in_1 ? 8'h41 : _GEN_1407; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1409 = 8'h81 == io_in_1 ? 8'h4f : _GEN_1408; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1410 = 8'h82 == io_in_1 ? 8'h5d : _GEN_1409; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1411 = 8'h83 == io_in_1 ? 8'h53 : _GEN_1410; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1412 = 8'h84 == io_in_1 ? 8'h79 : _GEN_1411; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1413 = 8'h85 == io_in_1 ? 8'h77 : _GEN_1412; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1414 = 8'h86 == io_in_1 ? 8'h65 : _GEN_1413; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1415 = 8'h87 == io_in_1 ? 8'h6b : _GEN_1414; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1416 = 8'h88 == io_in_1 ? 8'h31 : _GEN_1415; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1417 = 8'h89 == io_in_1 ? 8'h3f : _GEN_1416; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1418 = 8'h8a == io_in_1 ? 8'h2d : _GEN_1417; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1419 = 8'h8b == io_in_1 ? 8'h23 : _GEN_1418; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1420 = 8'h8c == io_in_1 ? 8'h9 : _GEN_1419; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1421 = 8'h8d == io_in_1 ? 8'h7 : _GEN_1420; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1422 = 8'h8e == io_in_1 ? 8'h15 : _GEN_1421; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1423 = 8'h8f == io_in_1 ? 8'h1b : _GEN_1422; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1424 = 8'h90 == io_in_1 ? 8'ha1 : _GEN_1423; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1425 = 8'h91 == io_in_1 ? 8'haf : _GEN_1424; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1426 = 8'h92 == io_in_1 ? 8'hbd : _GEN_1425; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1427 = 8'h93 == io_in_1 ? 8'hb3 : _GEN_1426; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1428 = 8'h94 == io_in_1 ? 8'h99 : _GEN_1427; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1429 = 8'h95 == io_in_1 ? 8'h97 : _GEN_1428; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1430 = 8'h96 == io_in_1 ? 8'h85 : _GEN_1429; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1431 = 8'h97 == io_in_1 ? 8'h8b : _GEN_1430; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1432 = 8'h98 == io_in_1 ? 8'hd1 : _GEN_1431; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1433 = 8'h99 == io_in_1 ? 8'hdf : _GEN_1432; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1434 = 8'h9a == io_in_1 ? 8'hcd : _GEN_1433; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1435 = 8'h9b == io_in_1 ? 8'hc3 : _GEN_1434; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1436 = 8'h9c == io_in_1 ? 8'he9 : _GEN_1435; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1437 = 8'h9d == io_in_1 ? 8'he7 : _GEN_1436; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1438 = 8'h9e == io_in_1 ? 8'hf5 : _GEN_1437; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1439 = 8'h9f == io_in_1 ? 8'hfb : _GEN_1438; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1440 = 8'ha0 == io_in_1 ? 8'h9a : _GEN_1439; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1441 = 8'ha1 == io_in_1 ? 8'h94 : _GEN_1440; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1442 = 8'ha2 == io_in_1 ? 8'h86 : _GEN_1441; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1443 = 8'ha3 == io_in_1 ? 8'h88 : _GEN_1442; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1444 = 8'ha4 == io_in_1 ? 8'ha2 : _GEN_1443; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1445 = 8'ha5 == io_in_1 ? 8'hac : _GEN_1444; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1446 = 8'ha6 == io_in_1 ? 8'hbe : _GEN_1445; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1447 = 8'ha7 == io_in_1 ? 8'hb0 : _GEN_1446; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1448 = 8'ha8 == io_in_1 ? 8'hea : _GEN_1447; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1449 = 8'ha9 == io_in_1 ? 8'he4 : _GEN_1448; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1450 = 8'haa == io_in_1 ? 8'hf6 : _GEN_1449; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1451 = 8'hab == io_in_1 ? 8'hf8 : _GEN_1450; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1452 = 8'hac == io_in_1 ? 8'hd2 : _GEN_1451; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1453 = 8'had == io_in_1 ? 8'hdc : _GEN_1452; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1454 = 8'hae == io_in_1 ? 8'hce : _GEN_1453; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1455 = 8'haf == io_in_1 ? 8'hc0 : _GEN_1454; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1456 = 8'hb0 == io_in_1 ? 8'h7a : _GEN_1455; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1457 = 8'hb1 == io_in_1 ? 8'h74 : _GEN_1456; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1458 = 8'hb2 == io_in_1 ? 8'h66 : _GEN_1457; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1459 = 8'hb3 == io_in_1 ? 8'h68 : _GEN_1458; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1460 = 8'hb4 == io_in_1 ? 8'h42 : _GEN_1459; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1461 = 8'hb5 == io_in_1 ? 8'h4c : _GEN_1460; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1462 = 8'hb6 == io_in_1 ? 8'h5e : _GEN_1461; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1463 = 8'hb7 == io_in_1 ? 8'h50 : _GEN_1462; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1464 = 8'hb8 == io_in_1 ? 8'ha : _GEN_1463; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1465 = 8'hb9 == io_in_1 ? 8'h4 : _GEN_1464; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1466 = 8'hba == io_in_1 ? 8'h16 : _GEN_1465; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1467 = 8'hbb == io_in_1 ? 8'h18 : _GEN_1466; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1468 = 8'hbc == io_in_1 ? 8'h32 : _GEN_1467; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1469 = 8'hbd == io_in_1 ? 8'h3c : _GEN_1468; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1470 = 8'hbe == io_in_1 ? 8'h2e : _GEN_1469; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1471 = 8'hbf == io_in_1 ? 8'h20 : _GEN_1470; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1472 = 8'hc0 == io_in_1 ? 8'hec : _GEN_1471; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1473 = 8'hc1 == io_in_1 ? 8'he2 : _GEN_1472; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1474 = 8'hc2 == io_in_1 ? 8'hf0 : _GEN_1473; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1475 = 8'hc3 == io_in_1 ? 8'hfe : _GEN_1474; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1476 = 8'hc4 == io_in_1 ? 8'hd4 : _GEN_1475; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1477 = 8'hc5 == io_in_1 ? 8'hda : _GEN_1476; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1478 = 8'hc6 == io_in_1 ? 8'hc8 : _GEN_1477; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1479 = 8'hc7 == io_in_1 ? 8'hc6 : _GEN_1478; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1480 = 8'hc8 == io_in_1 ? 8'h9c : _GEN_1479; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1481 = 8'hc9 == io_in_1 ? 8'h92 : _GEN_1480; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1482 = 8'hca == io_in_1 ? 8'h80 : _GEN_1481; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1483 = 8'hcb == io_in_1 ? 8'h8e : _GEN_1482; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1484 = 8'hcc == io_in_1 ? 8'ha4 : _GEN_1483; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1485 = 8'hcd == io_in_1 ? 8'haa : _GEN_1484; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1486 = 8'hce == io_in_1 ? 8'hb8 : _GEN_1485; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1487 = 8'hcf == io_in_1 ? 8'hb6 : _GEN_1486; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1488 = 8'hd0 == io_in_1 ? 8'hc : _GEN_1487; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1489 = 8'hd1 == io_in_1 ? 8'h2 : _GEN_1488; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1490 = 8'hd2 == io_in_1 ? 8'h10 : _GEN_1489; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1491 = 8'hd3 == io_in_1 ? 8'h1e : _GEN_1490; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1492 = 8'hd4 == io_in_1 ? 8'h34 : _GEN_1491; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1493 = 8'hd5 == io_in_1 ? 8'h3a : _GEN_1492; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1494 = 8'hd6 == io_in_1 ? 8'h28 : _GEN_1493; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1495 = 8'hd7 == io_in_1 ? 8'h26 : _GEN_1494; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1496 = 8'hd8 == io_in_1 ? 8'h7c : _GEN_1495; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1497 = 8'hd9 == io_in_1 ? 8'h72 : _GEN_1496; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1498 = 8'hda == io_in_1 ? 8'h60 : _GEN_1497; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1499 = 8'hdb == io_in_1 ? 8'h6e : _GEN_1498; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1500 = 8'hdc == io_in_1 ? 8'h44 : _GEN_1499; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1501 = 8'hdd == io_in_1 ? 8'h4a : _GEN_1500; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1502 = 8'hde == io_in_1 ? 8'h58 : _GEN_1501; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1503 = 8'hdf == io_in_1 ? 8'h56 : _GEN_1502; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1504 = 8'he0 == io_in_1 ? 8'h37 : _GEN_1503; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1505 = 8'he1 == io_in_1 ? 8'h39 : _GEN_1504; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1506 = 8'he2 == io_in_1 ? 8'h2b : _GEN_1505; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1507 = 8'he3 == io_in_1 ? 8'h25 : _GEN_1506; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1508 = 8'he4 == io_in_1 ? 8'hf : _GEN_1507; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1509 = 8'he5 == io_in_1 ? 8'h1 : _GEN_1508; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1510 = 8'he6 == io_in_1 ? 8'h13 : _GEN_1509; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1511 = 8'he7 == io_in_1 ? 8'h1d : _GEN_1510; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1512 = 8'he8 == io_in_1 ? 8'h47 : _GEN_1511; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1513 = 8'he9 == io_in_1 ? 8'h49 : _GEN_1512; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1514 = 8'hea == io_in_1 ? 8'h5b : _GEN_1513; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1515 = 8'heb == io_in_1 ? 8'h55 : _GEN_1514; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1516 = 8'hec == io_in_1 ? 8'h7f : _GEN_1515; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1517 = 8'hed == io_in_1 ? 8'h71 : _GEN_1516; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1518 = 8'hee == io_in_1 ? 8'h63 : _GEN_1517; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1519 = 8'hef == io_in_1 ? 8'h6d : _GEN_1518; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1520 = 8'hf0 == io_in_1 ? 8'hd7 : _GEN_1519; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1521 = 8'hf1 == io_in_1 ? 8'hd9 : _GEN_1520; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1522 = 8'hf2 == io_in_1 ? 8'hcb : _GEN_1521; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1523 = 8'hf3 == io_in_1 ? 8'hc5 : _GEN_1522; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1524 = 8'hf4 == io_in_1 ? 8'hef : _GEN_1523; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1525 = 8'hf5 == io_in_1 ? 8'he1 : _GEN_1524; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1526 = 8'hf6 == io_in_1 ? 8'hf3 : _GEN_1525; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1527 = 8'hf7 == io_in_1 ? 8'hfd : _GEN_1526; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1528 = 8'hf8 == io_in_1 ? 8'ha7 : _GEN_1527; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1529 = 8'hf9 == io_in_1 ? 8'ha9 : _GEN_1528; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1530 = 8'hfa == io_in_1 ? 8'hbb : _GEN_1529; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1531 = 8'hfb == io_in_1 ? 8'hb5 : _GEN_1530; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1532 = 8'hfc == io_in_1 ? 8'h9f : _GEN_1531; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1533 = 8'hfd == io_in_1 ? 8'h91 : _GEN_1532; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1534 = 8'hfe == io_in_1 ? 8'h83 : _GEN_1533; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1535 = 8'hff == io_in_1 ? 8'h8d : _GEN_1534; // @[AES_PipelinedElasticBuffer.scala 592:31 AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _T_3 = _GEN_1279 ^ _GEN_1535; // @[AES_PipelinedElasticBuffer.scala 592:31]
  wire [7:0] _GEN_1537 = 8'h1 == io_in_2 ? 8'hb : 8'h0; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1538 = 8'h2 == io_in_2 ? 8'h16 : _GEN_1537; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1539 = 8'h3 == io_in_2 ? 8'h1d : _GEN_1538; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1540 = 8'h4 == io_in_2 ? 8'h2c : _GEN_1539; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1541 = 8'h5 == io_in_2 ? 8'h27 : _GEN_1540; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1542 = 8'h6 == io_in_2 ? 8'h3a : _GEN_1541; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1543 = 8'h7 == io_in_2 ? 8'h31 : _GEN_1542; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1544 = 8'h8 == io_in_2 ? 8'h58 : _GEN_1543; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1545 = 8'h9 == io_in_2 ? 8'h53 : _GEN_1544; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1546 = 8'ha == io_in_2 ? 8'h4e : _GEN_1545; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1547 = 8'hb == io_in_2 ? 8'h45 : _GEN_1546; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1548 = 8'hc == io_in_2 ? 8'h74 : _GEN_1547; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1549 = 8'hd == io_in_2 ? 8'h7f : _GEN_1548; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1550 = 8'he == io_in_2 ? 8'h62 : _GEN_1549; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1551 = 8'hf == io_in_2 ? 8'h69 : _GEN_1550; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1552 = 8'h10 == io_in_2 ? 8'hb0 : _GEN_1551; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1553 = 8'h11 == io_in_2 ? 8'hbb : _GEN_1552; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1554 = 8'h12 == io_in_2 ? 8'ha6 : _GEN_1553; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1555 = 8'h13 == io_in_2 ? 8'had : _GEN_1554; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1556 = 8'h14 == io_in_2 ? 8'h9c : _GEN_1555; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1557 = 8'h15 == io_in_2 ? 8'h97 : _GEN_1556; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1558 = 8'h16 == io_in_2 ? 8'h8a : _GEN_1557; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1559 = 8'h17 == io_in_2 ? 8'h81 : _GEN_1558; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1560 = 8'h18 == io_in_2 ? 8'he8 : _GEN_1559; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1561 = 8'h19 == io_in_2 ? 8'he3 : _GEN_1560; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1562 = 8'h1a == io_in_2 ? 8'hfe : _GEN_1561; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1563 = 8'h1b == io_in_2 ? 8'hf5 : _GEN_1562; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1564 = 8'h1c == io_in_2 ? 8'hc4 : _GEN_1563; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1565 = 8'h1d == io_in_2 ? 8'hcf : _GEN_1564; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1566 = 8'h1e == io_in_2 ? 8'hd2 : _GEN_1565; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1567 = 8'h1f == io_in_2 ? 8'hd9 : _GEN_1566; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1568 = 8'h20 == io_in_2 ? 8'h7b : _GEN_1567; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1569 = 8'h21 == io_in_2 ? 8'h70 : _GEN_1568; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1570 = 8'h22 == io_in_2 ? 8'h6d : _GEN_1569; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1571 = 8'h23 == io_in_2 ? 8'h66 : _GEN_1570; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1572 = 8'h24 == io_in_2 ? 8'h57 : _GEN_1571; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1573 = 8'h25 == io_in_2 ? 8'h5c : _GEN_1572; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1574 = 8'h26 == io_in_2 ? 8'h41 : _GEN_1573; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1575 = 8'h27 == io_in_2 ? 8'h4a : _GEN_1574; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1576 = 8'h28 == io_in_2 ? 8'h23 : _GEN_1575; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1577 = 8'h29 == io_in_2 ? 8'h28 : _GEN_1576; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1578 = 8'h2a == io_in_2 ? 8'h35 : _GEN_1577; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1579 = 8'h2b == io_in_2 ? 8'h3e : _GEN_1578; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1580 = 8'h2c == io_in_2 ? 8'hf : _GEN_1579; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1581 = 8'h2d == io_in_2 ? 8'h4 : _GEN_1580; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1582 = 8'h2e == io_in_2 ? 8'h19 : _GEN_1581; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1583 = 8'h2f == io_in_2 ? 8'h12 : _GEN_1582; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1584 = 8'h30 == io_in_2 ? 8'hcb : _GEN_1583; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1585 = 8'h31 == io_in_2 ? 8'hc0 : _GEN_1584; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1586 = 8'h32 == io_in_2 ? 8'hdd : _GEN_1585; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1587 = 8'h33 == io_in_2 ? 8'hd6 : _GEN_1586; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1588 = 8'h34 == io_in_2 ? 8'he7 : _GEN_1587; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1589 = 8'h35 == io_in_2 ? 8'hec : _GEN_1588; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1590 = 8'h36 == io_in_2 ? 8'hf1 : _GEN_1589; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1591 = 8'h37 == io_in_2 ? 8'hfa : _GEN_1590; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1592 = 8'h38 == io_in_2 ? 8'h93 : _GEN_1591; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1593 = 8'h39 == io_in_2 ? 8'h98 : _GEN_1592; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1594 = 8'h3a == io_in_2 ? 8'h85 : _GEN_1593; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1595 = 8'h3b == io_in_2 ? 8'h8e : _GEN_1594; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1596 = 8'h3c == io_in_2 ? 8'hbf : _GEN_1595; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1597 = 8'h3d == io_in_2 ? 8'hb4 : _GEN_1596; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1598 = 8'h3e == io_in_2 ? 8'ha9 : _GEN_1597; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1599 = 8'h3f == io_in_2 ? 8'ha2 : _GEN_1598; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1600 = 8'h40 == io_in_2 ? 8'hf6 : _GEN_1599; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1601 = 8'h41 == io_in_2 ? 8'hfd : _GEN_1600; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1602 = 8'h42 == io_in_2 ? 8'he0 : _GEN_1601; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1603 = 8'h43 == io_in_2 ? 8'heb : _GEN_1602; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1604 = 8'h44 == io_in_2 ? 8'hda : _GEN_1603; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1605 = 8'h45 == io_in_2 ? 8'hd1 : _GEN_1604; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1606 = 8'h46 == io_in_2 ? 8'hcc : _GEN_1605; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1607 = 8'h47 == io_in_2 ? 8'hc7 : _GEN_1606; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1608 = 8'h48 == io_in_2 ? 8'hae : _GEN_1607; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1609 = 8'h49 == io_in_2 ? 8'ha5 : _GEN_1608; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1610 = 8'h4a == io_in_2 ? 8'hb8 : _GEN_1609; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1611 = 8'h4b == io_in_2 ? 8'hb3 : _GEN_1610; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1612 = 8'h4c == io_in_2 ? 8'h82 : _GEN_1611; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1613 = 8'h4d == io_in_2 ? 8'h89 : _GEN_1612; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1614 = 8'h4e == io_in_2 ? 8'h94 : _GEN_1613; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1615 = 8'h4f == io_in_2 ? 8'h9f : _GEN_1614; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1616 = 8'h50 == io_in_2 ? 8'h46 : _GEN_1615; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1617 = 8'h51 == io_in_2 ? 8'h4d : _GEN_1616; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1618 = 8'h52 == io_in_2 ? 8'h50 : _GEN_1617; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1619 = 8'h53 == io_in_2 ? 8'h5b : _GEN_1618; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1620 = 8'h54 == io_in_2 ? 8'h6a : _GEN_1619; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1621 = 8'h55 == io_in_2 ? 8'h61 : _GEN_1620; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1622 = 8'h56 == io_in_2 ? 8'h7c : _GEN_1621; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1623 = 8'h57 == io_in_2 ? 8'h77 : _GEN_1622; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1624 = 8'h58 == io_in_2 ? 8'h1e : _GEN_1623; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1625 = 8'h59 == io_in_2 ? 8'h15 : _GEN_1624; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1626 = 8'h5a == io_in_2 ? 8'h8 : _GEN_1625; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1627 = 8'h5b == io_in_2 ? 8'h3 : _GEN_1626; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1628 = 8'h5c == io_in_2 ? 8'h32 : _GEN_1627; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1629 = 8'h5d == io_in_2 ? 8'h39 : _GEN_1628; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1630 = 8'h5e == io_in_2 ? 8'h24 : _GEN_1629; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1631 = 8'h5f == io_in_2 ? 8'h2f : _GEN_1630; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1632 = 8'h60 == io_in_2 ? 8'h8d : _GEN_1631; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1633 = 8'h61 == io_in_2 ? 8'h86 : _GEN_1632; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1634 = 8'h62 == io_in_2 ? 8'h9b : _GEN_1633; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1635 = 8'h63 == io_in_2 ? 8'h90 : _GEN_1634; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1636 = 8'h64 == io_in_2 ? 8'ha1 : _GEN_1635; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1637 = 8'h65 == io_in_2 ? 8'haa : _GEN_1636; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1638 = 8'h66 == io_in_2 ? 8'hb7 : _GEN_1637; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1639 = 8'h67 == io_in_2 ? 8'hbc : _GEN_1638; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1640 = 8'h68 == io_in_2 ? 8'hd5 : _GEN_1639; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1641 = 8'h69 == io_in_2 ? 8'hde : _GEN_1640; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1642 = 8'h6a == io_in_2 ? 8'hc3 : _GEN_1641; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1643 = 8'h6b == io_in_2 ? 8'hc8 : _GEN_1642; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1644 = 8'h6c == io_in_2 ? 8'hf9 : _GEN_1643; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1645 = 8'h6d == io_in_2 ? 8'hf2 : _GEN_1644; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1646 = 8'h6e == io_in_2 ? 8'hef : _GEN_1645; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1647 = 8'h6f == io_in_2 ? 8'he4 : _GEN_1646; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1648 = 8'h70 == io_in_2 ? 8'h3d : _GEN_1647; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1649 = 8'h71 == io_in_2 ? 8'h36 : _GEN_1648; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1650 = 8'h72 == io_in_2 ? 8'h2b : _GEN_1649; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1651 = 8'h73 == io_in_2 ? 8'h20 : _GEN_1650; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1652 = 8'h74 == io_in_2 ? 8'h11 : _GEN_1651; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1653 = 8'h75 == io_in_2 ? 8'h1a : _GEN_1652; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1654 = 8'h76 == io_in_2 ? 8'h7 : _GEN_1653; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1655 = 8'h77 == io_in_2 ? 8'hc : _GEN_1654; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1656 = 8'h78 == io_in_2 ? 8'h65 : _GEN_1655; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1657 = 8'h79 == io_in_2 ? 8'h6e : _GEN_1656; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1658 = 8'h7a == io_in_2 ? 8'h73 : _GEN_1657; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1659 = 8'h7b == io_in_2 ? 8'h78 : _GEN_1658; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1660 = 8'h7c == io_in_2 ? 8'h49 : _GEN_1659; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1661 = 8'h7d == io_in_2 ? 8'h42 : _GEN_1660; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1662 = 8'h7e == io_in_2 ? 8'h5f : _GEN_1661; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1663 = 8'h7f == io_in_2 ? 8'h54 : _GEN_1662; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1664 = 8'h80 == io_in_2 ? 8'hf7 : _GEN_1663; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1665 = 8'h81 == io_in_2 ? 8'hfc : _GEN_1664; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1666 = 8'h82 == io_in_2 ? 8'he1 : _GEN_1665; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1667 = 8'h83 == io_in_2 ? 8'hea : _GEN_1666; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1668 = 8'h84 == io_in_2 ? 8'hdb : _GEN_1667; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1669 = 8'h85 == io_in_2 ? 8'hd0 : _GEN_1668; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1670 = 8'h86 == io_in_2 ? 8'hcd : _GEN_1669; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1671 = 8'h87 == io_in_2 ? 8'hc6 : _GEN_1670; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1672 = 8'h88 == io_in_2 ? 8'haf : _GEN_1671; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1673 = 8'h89 == io_in_2 ? 8'ha4 : _GEN_1672; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1674 = 8'h8a == io_in_2 ? 8'hb9 : _GEN_1673; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1675 = 8'h8b == io_in_2 ? 8'hb2 : _GEN_1674; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1676 = 8'h8c == io_in_2 ? 8'h83 : _GEN_1675; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1677 = 8'h8d == io_in_2 ? 8'h88 : _GEN_1676; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1678 = 8'h8e == io_in_2 ? 8'h95 : _GEN_1677; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1679 = 8'h8f == io_in_2 ? 8'h9e : _GEN_1678; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1680 = 8'h90 == io_in_2 ? 8'h47 : _GEN_1679; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1681 = 8'h91 == io_in_2 ? 8'h4c : _GEN_1680; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1682 = 8'h92 == io_in_2 ? 8'h51 : _GEN_1681; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1683 = 8'h93 == io_in_2 ? 8'h5a : _GEN_1682; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1684 = 8'h94 == io_in_2 ? 8'h6b : _GEN_1683; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1685 = 8'h95 == io_in_2 ? 8'h60 : _GEN_1684; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1686 = 8'h96 == io_in_2 ? 8'h7d : _GEN_1685; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1687 = 8'h97 == io_in_2 ? 8'h76 : _GEN_1686; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1688 = 8'h98 == io_in_2 ? 8'h1f : _GEN_1687; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1689 = 8'h99 == io_in_2 ? 8'h14 : _GEN_1688; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1690 = 8'h9a == io_in_2 ? 8'h9 : _GEN_1689; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1691 = 8'h9b == io_in_2 ? 8'h2 : _GEN_1690; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1692 = 8'h9c == io_in_2 ? 8'h33 : _GEN_1691; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1693 = 8'h9d == io_in_2 ? 8'h38 : _GEN_1692; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1694 = 8'h9e == io_in_2 ? 8'h25 : _GEN_1693; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1695 = 8'h9f == io_in_2 ? 8'h2e : _GEN_1694; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1696 = 8'ha0 == io_in_2 ? 8'h8c : _GEN_1695; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1697 = 8'ha1 == io_in_2 ? 8'h87 : _GEN_1696; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1698 = 8'ha2 == io_in_2 ? 8'h9a : _GEN_1697; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1699 = 8'ha3 == io_in_2 ? 8'h91 : _GEN_1698; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1700 = 8'ha4 == io_in_2 ? 8'ha0 : _GEN_1699; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1701 = 8'ha5 == io_in_2 ? 8'hab : _GEN_1700; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1702 = 8'ha6 == io_in_2 ? 8'hb6 : _GEN_1701; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1703 = 8'ha7 == io_in_2 ? 8'hbd : _GEN_1702; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1704 = 8'ha8 == io_in_2 ? 8'hd4 : _GEN_1703; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1705 = 8'ha9 == io_in_2 ? 8'hdf : _GEN_1704; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1706 = 8'haa == io_in_2 ? 8'hc2 : _GEN_1705; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1707 = 8'hab == io_in_2 ? 8'hc9 : _GEN_1706; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1708 = 8'hac == io_in_2 ? 8'hf8 : _GEN_1707; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1709 = 8'had == io_in_2 ? 8'hf3 : _GEN_1708; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1710 = 8'hae == io_in_2 ? 8'hee : _GEN_1709; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1711 = 8'haf == io_in_2 ? 8'he5 : _GEN_1710; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1712 = 8'hb0 == io_in_2 ? 8'h3c : _GEN_1711; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1713 = 8'hb1 == io_in_2 ? 8'h37 : _GEN_1712; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1714 = 8'hb2 == io_in_2 ? 8'h2a : _GEN_1713; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1715 = 8'hb3 == io_in_2 ? 8'h21 : _GEN_1714; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1716 = 8'hb4 == io_in_2 ? 8'h10 : _GEN_1715; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1717 = 8'hb5 == io_in_2 ? 8'h1b : _GEN_1716; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1718 = 8'hb6 == io_in_2 ? 8'h6 : _GEN_1717; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1719 = 8'hb7 == io_in_2 ? 8'hd : _GEN_1718; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1720 = 8'hb8 == io_in_2 ? 8'h64 : _GEN_1719; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1721 = 8'hb9 == io_in_2 ? 8'h6f : _GEN_1720; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1722 = 8'hba == io_in_2 ? 8'h72 : _GEN_1721; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1723 = 8'hbb == io_in_2 ? 8'h79 : _GEN_1722; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1724 = 8'hbc == io_in_2 ? 8'h48 : _GEN_1723; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1725 = 8'hbd == io_in_2 ? 8'h43 : _GEN_1724; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1726 = 8'hbe == io_in_2 ? 8'h5e : _GEN_1725; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1727 = 8'hbf == io_in_2 ? 8'h55 : _GEN_1726; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1728 = 8'hc0 == io_in_2 ? 8'h1 : _GEN_1727; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1729 = 8'hc1 == io_in_2 ? 8'ha : _GEN_1728; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1730 = 8'hc2 == io_in_2 ? 8'h17 : _GEN_1729; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1731 = 8'hc3 == io_in_2 ? 8'h1c : _GEN_1730; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1732 = 8'hc4 == io_in_2 ? 8'h2d : _GEN_1731; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1733 = 8'hc5 == io_in_2 ? 8'h26 : _GEN_1732; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1734 = 8'hc6 == io_in_2 ? 8'h3b : _GEN_1733; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1735 = 8'hc7 == io_in_2 ? 8'h30 : _GEN_1734; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1736 = 8'hc8 == io_in_2 ? 8'h59 : _GEN_1735; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1737 = 8'hc9 == io_in_2 ? 8'h52 : _GEN_1736; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1738 = 8'hca == io_in_2 ? 8'h4f : _GEN_1737; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1739 = 8'hcb == io_in_2 ? 8'h44 : _GEN_1738; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1740 = 8'hcc == io_in_2 ? 8'h75 : _GEN_1739; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1741 = 8'hcd == io_in_2 ? 8'h7e : _GEN_1740; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1742 = 8'hce == io_in_2 ? 8'h63 : _GEN_1741; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1743 = 8'hcf == io_in_2 ? 8'h68 : _GEN_1742; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1744 = 8'hd0 == io_in_2 ? 8'hb1 : _GEN_1743; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1745 = 8'hd1 == io_in_2 ? 8'hba : _GEN_1744; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1746 = 8'hd2 == io_in_2 ? 8'ha7 : _GEN_1745; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1747 = 8'hd3 == io_in_2 ? 8'hac : _GEN_1746; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1748 = 8'hd4 == io_in_2 ? 8'h9d : _GEN_1747; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1749 = 8'hd5 == io_in_2 ? 8'h96 : _GEN_1748; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1750 = 8'hd6 == io_in_2 ? 8'h8b : _GEN_1749; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1751 = 8'hd7 == io_in_2 ? 8'h80 : _GEN_1750; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1752 = 8'hd8 == io_in_2 ? 8'he9 : _GEN_1751; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1753 = 8'hd9 == io_in_2 ? 8'he2 : _GEN_1752; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1754 = 8'hda == io_in_2 ? 8'hff : _GEN_1753; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1755 = 8'hdb == io_in_2 ? 8'hf4 : _GEN_1754; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1756 = 8'hdc == io_in_2 ? 8'hc5 : _GEN_1755; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1757 = 8'hdd == io_in_2 ? 8'hce : _GEN_1756; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1758 = 8'hde == io_in_2 ? 8'hd3 : _GEN_1757; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1759 = 8'hdf == io_in_2 ? 8'hd8 : _GEN_1758; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1760 = 8'he0 == io_in_2 ? 8'h7a : _GEN_1759; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1761 = 8'he1 == io_in_2 ? 8'h71 : _GEN_1760; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1762 = 8'he2 == io_in_2 ? 8'h6c : _GEN_1761; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1763 = 8'he3 == io_in_2 ? 8'h67 : _GEN_1762; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1764 = 8'he4 == io_in_2 ? 8'h56 : _GEN_1763; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1765 = 8'he5 == io_in_2 ? 8'h5d : _GEN_1764; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1766 = 8'he6 == io_in_2 ? 8'h40 : _GEN_1765; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1767 = 8'he7 == io_in_2 ? 8'h4b : _GEN_1766; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1768 = 8'he8 == io_in_2 ? 8'h22 : _GEN_1767; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1769 = 8'he9 == io_in_2 ? 8'h29 : _GEN_1768; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1770 = 8'hea == io_in_2 ? 8'h34 : _GEN_1769; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1771 = 8'heb == io_in_2 ? 8'h3f : _GEN_1770; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1772 = 8'hec == io_in_2 ? 8'he : _GEN_1771; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1773 = 8'hed == io_in_2 ? 8'h5 : _GEN_1772; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1774 = 8'hee == io_in_2 ? 8'h18 : _GEN_1773; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1775 = 8'hef == io_in_2 ? 8'h13 : _GEN_1774; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1776 = 8'hf0 == io_in_2 ? 8'hca : _GEN_1775; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1777 = 8'hf1 == io_in_2 ? 8'hc1 : _GEN_1776; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1778 = 8'hf2 == io_in_2 ? 8'hdc : _GEN_1777; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1779 = 8'hf3 == io_in_2 ? 8'hd7 : _GEN_1778; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1780 = 8'hf4 == io_in_2 ? 8'he6 : _GEN_1779; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1781 = 8'hf5 == io_in_2 ? 8'hed : _GEN_1780; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1782 = 8'hf6 == io_in_2 ? 8'hf0 : _GEN_1781; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1783 = 8'hf7 == io_in_2 ? 8'hfb : _GEN_1782; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1784 = 8'hf8 == io_in_2 ? 8'h92 : _GEN_1783; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1785 = 8'hf9 == io_in_2 ? 8'h99 : _GEN_1784; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1786 = 8'hfa == io_in_2 ? 8'h84 : _GEN_1785; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1787 = 8'hfb == io_in_2 ? 8'h8f : _GEN_1786; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1788 = 8'hfc == io_in_2 ? 8'hbe : _GEN_1787; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1789 = 8'hfd == io_in_2 ? 8'hb5 : _GEN_1788; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1790 = 8'hfe == io_in_2 ? 8'ha8 : _GEN_1789; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1791 = 8'hff == io_in_2 ? 8'ha3 : _GEN_1790; // @[AES_PipelinedElasticBuffer.scala 592:49 AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _T_4 = _T_3 ^ _GEN_1791; // @[AES_PipelinedElasticBuffer.scala 592:49]
  wire [7:0] _GEN_1793 = 8'h1 == io_in_3 ? 8'hd : 8'h0; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1794 = 8'h2 == io_in_3 ? 8'h1a : _GEN_1793; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1795 = 8'h3 == io_in_3 ? 8'h17 : _GEN_1794; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1796 = 8'h4 == io_in_3 ? 8'h34 : _GEN_1795; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1797 = 8'h5 == io_in_3 ? 8'h39 : _GEN_1796; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1798 = 8'h6 == io_in_3 ? 8'h2e : _GEN_1797; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1799 = 8'h7 == io_in_3 ? 8'h23 : _GEN_1798; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1800 = 8'h8 == io_in_3 ? 8'h68 : _GEN_1799; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1801 = 8'h9 == io_in_3 ? 8'h65 : _GEN_1800; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1802 = 8'ha == io_in_3 ? 8'h72 : _GEN_1801; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1803 = 8'hb == io_in_3 ? 8'h7f : _GEN_1802; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1804 = 8'hc == io_in_3 ? 8'h5c : _GEN_1803; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1805 = 8'hd == io_in_3 ? 8'h51 : _GEN_1804; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1806 = 8'he == io_in_3 ? 8'h46 : _GEN_1805; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1807 = 8'hf == io_in_3 ? 8'h4b : _GEN_1806; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1808 = 8'h10 == io_in_3 ? 8'hd0 : _GEN_1807; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1809 = 8'h11 == io_in_3 ? 8'hdd : _GEN_1808; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1810 = 8'h12 == io_in_3 ? 8'hca : _GEN_1809; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1811 = 8'h13 == io_in_3 ? 8'hc7 : _GEN_1810; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1812 = 8'h14 == io_in_3 ? 8'he4 : _GEN_1811; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1813 = 8'h15 == io_in_3 ? 8'he9 : _GEN_1812; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1814 = 8'h16 == io_in_3 ? 8'hfe : _GEN_1813; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1815 = 8'h17 == io_in_3 ? 8'hf3 : _GEN_1814; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1816 = 8'h18 == io_in_3 ? 8'hb8 : _GEN_1815; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1817 = 8'h19 == io_in_3 ? 8'hb5 : _GEN_1816; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1818 = 8'h1a == io_in_3 ? 8'ha2 : _GEN_1817; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1819 = 8'h1b == io_in_3 ? 8'haf : _GEN_1818; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1820 = 8'h1c == io_in_3 ? 8'h8c : _GEN_1819; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1821 = 8'h1d == io_in_3 ? 8'h81 : _GEN_1820; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1822 = 8'h1e == io_in_3 ? 8'h96 : _GEN_1821; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1823 = 8'h1f == io_in_3 ? 8'h9b : _GEN_1822; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1824 = 8'h20 == io_in_3 ? 8'hbb : _GEN_1823; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1825 = 8'h21 == io_in_3 ? 8'hb6 : _GEN_1824; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1826 = 8'h22 == io_in_3 ? 8'ha1 : _GEN_1825; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1827 = 8'h23 == io_in_3 ? 8'hac : _GEN_1826; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1828 = 8'h24 == io_in_3 ? 8'h8f : _GEN_1827; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1829 = 8'h25 == io_in_3 ? 8'h82 : _GEN_1828; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1830 = 8'h26 == io_in_3 ? 8'h95 : _GEN_1829; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1831 = 8'h27 == io_in_3 ? 8'h98 : _GEN_1830; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1832 = 8'h28 == io_in_3 ? 8'hd3 : _GEN_1831; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1833 = 8'h29 == io_in_3 ? 8'hde : _GEN_1832; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1834 = 8'h2a == io_in_3 ? 8'hc9 : _GEN_1833; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1835 = 8'h2b == io_in_3 ? 8'hc4 : _GEN_1834; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1836 = 8'h2c == io_in_3 ? 8'he7 : _GEN_1835; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1837 = 8'h2d == io_in_3 ? 8'hea : _GEN_1836; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1838 = 8'h2e == io_in_3 ? 8'hfd : _GEN_1837; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1839 = 8'h2f == io_in_3 ? 8'hf0 : _GEN_1838; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1840 = 8'h30 == io_in_3 ? 8'h6b : _GEN_1839; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1841 = 8'h31 == io_in_3 ? 8'h66 : _GEN_1840; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1842 = 8'h32 == io_in_3 ? 8'h71 : _GEN_1841; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1843 = 8'h33 == io_in_3 ? 8'h7c : _GEN_1842; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1844 = 8'h34 == io_in_3 ? 8'h5f : _GEN_1843; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1845 = 8'h35 == io_in_3 ? 8'h52 : _GEN_1844; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1846 = 8'h36 == io_in_3 ? 8'h45 : _GEN_1845; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1847 = 8'h37 == io_in_3 ? 8'h48 : _GEN_1846; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1848 = 8'h38 == io_in_3 ? 8'h3 : _GEN_1847; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1849 = 8'h39 == io_in_3 ? 8'he : _GEN_1848; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1850 = 8'h3a == io_in_3 ? 8'h19 : _GEN_1849; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1851 = 8'h3b == io_in_3 ? 8'h14 : _GEN_1850; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1852 = 8'h3c == io_in_3 ? 8'h37 : _GEN_1851; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1853 = 8'h3d == io_in_3 ? 8'h3a : _GEN_1852; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1854 = 8'h3e == io_in_3 ? 8'h2d : _GEN_1853; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1855 = 8'h3f == io_in_3 ? 8'h20 : _GEN_1854; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1856 = 8'h40 == io_in_3 ? 8'h6d : _GEN_1855; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1857 = 8'h41 == io_in_3 ? 8'h60 : _GEN_1856; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1858 = 8'h42 == io_in_3 ? 8'h77 : _GEN_1857; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1859 = 8'h43 == io_in_3 ? 8'h7a : _GEN_1858; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1860 = 8'h44 == io_in_3 ? 8'h59 : _GEN_1859; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1861 = 8'h45 == io_in_3 ? 8'h54 : _GEN_1860; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1862 = 8'h46 == io_in_3 ? 8'h43 : _GEN_1861; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1863 = 8'h47 == io_in_3 ? 8'h4e : _GEN_1862; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1864 = 8'h48 == io_in_3 ? 8'h5 : _GEN_1863; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1865 = 8'h49 == io_in_3 ? 8'h8 : _GEN_1864; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1866 = 8'h4a == io_in_3 ? 8'h1f : _GEN_1865; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1867 = 8'h4b == io_in_3 ? 8'h12 : _GEN_1866; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1868 = 8'h4c == io_in_3 ? 8'h31 : _GEN_1867; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1869 = 8'h4d == io_in_3 ? 8'h3c : _GEN_1868; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1870 = 8'h4e == io_in_3 ? 8'h2b : _GEN_1869; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1871 = 8'h4f == io_in_3 ? 8'h26 : _GEN_1870; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1872 = 8'h50 == io_in_3 ? 8'hbd : _GEN_1871; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1873 = 8'h51 == io_in_3 ? 8'hb0 : _GEN_1872; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1874 = 8'h52 == io_in_3 ? 8'ha7 : _GEN_1873; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1875 = 8'h53 == io_in_3 ? 8'haa : _GEN_1874; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1876 = 8'h54 == io_in_3 ? 8'h89 : _GEN_1875; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1877 = 8'h55 == io_in_3 ? 8'h84 : _GEN_1876; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1878 = 8'h56 == io_in_3 ? 8'h93 : _GEN_1877; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1879 = 8'h57 == io_in_3 ? 8'h9e : _GEN_1878; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1880 = 8'h58 == io_in_3 ? 8'hd5 : _GEN_1879; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1881 = 8'h59 == io_in_3 ? 8'hd8 : _GEN_1880; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1882 = 8'h5a == io_in_3 ? 8'hcf : _GEN_1881; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1883 = 8'h5b == io_in_3 ? 8'hc2 : _GEN_1882; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1884 = 8'h5c == io_in_3 ? 8'he1 : _GEN_1883; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1885 = 8'h5d == io_in_3 ? 8'hec : _GEN_1884; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1886 = 8'h5e == io_in_3 ? 8'hfb : _GEN_1885; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1887 = 8'h5f == io_in_3 ? 8'hf6 : _GEN_1886; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1888 = 8'h60 == io_in_3 ? 8'hd6 : _GEN_1887; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1889 = 8'h61 == io_in_3 ? 8'hdb : _GEN_1888; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1890 = 8'h62 == io_in_3 ? 8'hcc : _GEN_1889; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1891 = 8'h63 == io_in_3 ? 8'hc1 : _GEN_1890; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1892 = 8'h64 == io_in_3 ? 8'he2 : _GEN_1891; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1893 = 8'h65 == io_in_3 ? 8'hef : _GEN_1892; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1894 = 8'h66 == io_in_3 ? 8'hf8 : _GEN_1893; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1895 = 8'h67 == io_in_3 ? 8'hf5 : _GEN_1894; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1896 = 8'h68 == io_in_3 ? 8'hbe : _GEN_1895; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1897 = 8'h69 == io_in_3 ? 8'hb3 : _GEN_1896; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1898 = 8'h6a == io_in_3 ? 8'ha4 : _GEN_1897; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1899 = 8'h6b == io_in_3 ? 8'ha9 : _GEN_1898; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1900 = 8'h6c == io_in_3 ? 8'h8a : _GEN_1899; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1901 = 8'h6d == io_in_3 ? 8'h87 : _GEN_1900; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1902 = 8'h6e == io_in_3 ? 8'h90 : _GEN_1901; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1903 = 8'h6f == io_in_3 ? 8'h9d : _GEN_1902; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1904 = 8'h70 == io_in_3 ? 8'h6 : _GEN_1903; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1905 = 8'h71 == io_in_3 ? 8'hb : _GEN_1904; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1906 = 8'h72 == io_in_3 ? 8'h1c : _GEN_1905; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1907 = 8'h73 == io_in_3 ? 8'h11 : _GEN_1906; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1908 = 8'h74 == io_in_3 ? 8'h32 : _GEN_1907; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1909 = 8'h75 == io_in_3 ? 8'h3f : _GEN_1908; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1910 = 8'h76 == io_in_3 ? 8'h28 : _GEN_1909; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1911 = 8'h77 == io_in_3 ? 8'h25 : _GEN_1910; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1912 = 8'h78 == io_in_3 ? 8'h6e : _GEN_1911; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1913 = 8'h79 == io_in_3 ? 8'h63 : _GEN_1912; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1914 = 8'h7a == io_in_3 ? 8'h74 : _GEN_1913; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1915 = 8'h7b == io_in_3 ? 8'h79 : _GEN_1914; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1916 = 8'h7c == io_in_3 ? 8'h5a : _GEN_1915; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1917 = 8'h7d == io_in_3 ? 8'h57 : _GEN_1916; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1918 = 8'h7e == io_in_3 ? 8'h40 : _GEN_1917; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1919 = 8'h7f == io_in_3 ? 8'h4d : _GEN_1918; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1920 = 8'h80 == io_in_3 ? 8'hda : _GEN_1919; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1921 = 8'h81 == io_in_3 ? 8'hd7 : _GEN_1920; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1922 = 8'h82 == io_in_3 ? 8'hc0 : _GEN_1921; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1923 = 8'h83 == io_in_3 ? 8'hcd : _GEN_1922; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1924 = 8'h84 == io_in_3 ? 8'hee : _GEN_1923; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1925 = 8'h85 == io_in_3 ? 8'he3 : _GEN_1924; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1926 = 8'h86 == io_in_3 ? 8'hf4 : _GEN_1925; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1927 = 8'h87 == io_in_3 ? 8'hf9 : _GEN_1926; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1928 = 8'h88 == io_in_3 ? 8'hb2 : _GEN_1927; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1929 = 8'h89 == io_in_3 ? 8'hbf : _GEN_1928; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1930 = 8'h8a == io_in_3 ? 8'ha8 : _GEN_1929; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1931 = 8'h8b == io_in_3 ? 8'ha5 : _GEN_1930; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1932 = 8'h8c == io_in_3 ? 8'h86 : _GEN_1931; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1933 = 8'h8d == io_in_3 ? 8'h8b : _GEN_1932; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1934 = 8'h8e == io_in_3 ? 8'h9c : _GEN_1933; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1935 = 8'h8f == io_in_3 ? 8'h91 : _GEN_1934; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1936 = 8'h90 == io_in_3 ? 8'ha : _GEN_1935; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1937 = 8'h91 == io_in_3 ? 8'h7 : _GEN_1936; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1938 = 8'h92 == io_in_3 ? 8'h10 : _GEN_1937; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1939 = 8'h93 == io_in_3 ? 8'h1d : _GEN_1938; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1940 = 8'h94 == io_in_3 ? 8'h3e : _GEN_1939; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1941 = 8'h95 == io_in_3 ? 8'h33 : _GEN_1940; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1942 = 8'h96 == io_in_3 ? 8'h24 : _GEN_1941; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1943 = 8'h97 == io_in_3 ? 8'h29 : _GEN_1942; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1944 = 8'h98 == io_in_3 ? 8'h62 : _GEN_1943; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1945 = 8'h99 == io_in_3 ? 8'h6f : _GEN_1944; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1946 = 8'h9a == io_in_3 ? 8'h78 : _GEN_1945; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1947 = 8'h9b == io_in_3 ? 8'h75 : _GEN_1946; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1948 = 8'h9c == io_in_3 ? 8'h56 : _GEN_1947; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1949 = 8'h9d == io_in_3 ? 8'h5b : _GEN_1948; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1950 = 8'h9e == io_in_3 ? 8'h4c : _GEN_1949; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1951 = 8'h9f == io_in_3 ? 8'h41 : _GEN_1950; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1952 = 8'ha0 == io_in_3 ? 8'h61 : _GEN_1951; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1953 = 8'ha1 == io_in_3 ? 8'h6c : _GEN_1952; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1954 = 8'ha2 == io_in_3 ? 8'h7b : _GEN_1953; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1955 = 8'ha3 == io_in_3 ? 8'h76 : _GEN_1954; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1956 = 8'ha4 == io_in_3 ? 8'h55 : _GEN_1955; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1957 = 8'ha5 == io_in_3 ? 8'h58 : _GEN_1956; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1958 = 8'ha6 == io_in_3 ? 8'h4f : _GEN_1957; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1959 = 8'ha7 == io_in_3 ? 8'h42 : _GEN_1958; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1960 = 8'ha8 == io_in_3 ? 8'h9 : _GEN_1959; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1961 = 8'ha9 == io_in_3 ? 8'h4 : _GEN_1960; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1962 = 8'haa == io_in_3 ? 8'h13 : _GEN_1961; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1963 = 8'hab == io_in_3 ? 8'h1e : _GEN_1962; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1964 = 8'hac == io_in_3 ? 8'h3d : _GEN_1963; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1965 = 8'had == io_in_3 ? 8'h30 : _GEN_1964; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1966 = 8'hae == io_in_3 ? 8'h27 : _GEN_1965; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1967 = 8'haf == io_in_3 ? 8'h2a : _GEN_1966; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1968 = 8'hb0 == io_in_3 ? 8'hb1 : _GEN_1967; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1969 = 8'hb1 == io_in_3 ? 8'hbc : _GEN_1968; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1970 = 8'hb2 == io_in_3 ? 8'hab : _GEN_1969; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1971 = 8'hb3 == io_in_3 ? 8'ha6 : _GEN_1970; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1972 = 8'hb4 == io_in_3 ? 8'h85 : _GEN_1971; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1973 = 8'hb5 == io_in_3 ? 8'h88 : _GEN_1972; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1974 = 8'hb6 == io_in_3 ? 8'h9f : _GEN_1973; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1975 = 8'hb7 == io_in_3 ? 8'h92 : _GEN_1974; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1976 = 8'hb8 == io_in_3 ? 8'hd9 : _GEN_1975; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1977 = 8'hb9 == io_in_3 ? 8'hd4 : _GEN_1976; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1978 = 8'hba == io_in_3 ? 8'hc3 : _GEN_1977; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1979 = 8'hbb == io_in_3 ? 8'hce : _GEN_1978; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1980 = 8'hbc == io_in_3 ? 8'hed : _GEN_1979; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1981 = 8'hbd == io_in_3 ? 8'he0 : _GEN_1980; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1982 = 8'hbe == io_in_3 ? 8'hf7 : _GEN_1981; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1983 = 8'hbf == io_in_3 ? 8'hfa : _GEN_1982; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1984 = 8'hc0 == io_in_3 ? 8'hb7 : _GEN_1983; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1985 = 8'hc1 == io_in_3 ? 8'hba : _GEN_1984; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1986 = 8'hc2 == io_in_3 ? 8'had : _GEN_1985; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1987 = 8'hc3 == io_in_3 ? 8'ha0 : _GEN_1986; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1988 = 8'hc4 == io_in_3 ? 8'h83 : _GEN_1987; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1989 = 8'hc5 == io_in_3 ? 8'h8e : _GEN_1988; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1990 = 8'hc6 == io_in_3 ? 8'h99 : _GEN_1989; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1991 = 8'hc7 == io_in_3 ? 8'h94 : _GEN_1990; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1992 = 8'hc8 == io_in_3 ? 8'hdf : _GEN_1991; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1993 = 8'hc9 == io_in_3 ? 8'hd2 : _GEN_1992; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1994 = 8'hca == io_in_3 ? 8'hc5 : _GEN_1993; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1995 = 8'hcb == io_in_3 ? 8'hc8 : _GEN_1994; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1996 = 8'hcc == io_in_3 ? 8'heb : _GEN_1995; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1997 = 8'hcd == io_in_3 ? 8'he6 : _GEN_1996; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1998 = 8'hce == io_in_3 ? 8'hf1 : _GEN_1997; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_1999 = 8'hcf == io_in_3 ? 8'hfc : _GEN_1998; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2000 = 8'hd0 == io_in_3 ? 8'h67 : _GEN_1999; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2001 = 8'hd1 == io_in_3 ? 8'h6a : _GEN_2000; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2002 = 8'hd2 == io_in_3 ? 8'h7d : _GEN_2001; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2003 = 8'hd3 == io_in_3 ? 8'h70 : _GEN_2002; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2004 = 8'hd4 == io_in_3 ? 8'h53 : _GEN_2003; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2005 = 8'hd5 == io_in_3 ? 8'h5e : _GEN_2004; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2006 = 8'hd6 == io_in_3 ? 8'h49 : _GEN_2005; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2007 = 8'hd7 == io_in_3 ? 8'h44 : _GEN_2006; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2008 = 8'hd8 == io_in_3 ? 8'hf : _GEN_2007; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2009 = 8'hd9 == io_in_3 ? 8'h2 : _GEN_2008; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2010 = 8'hda == io_in_3 ? 8'h15 : _GEN_2009; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2011 = 8'hdb == io_in_3 ? 8'h18 : _GEN_2010; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2012 = 8'hdc == io_in_3 ? 8'h3b : _GEN_2011; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2013 = 8'hdd == io_in_3 ? 8'h36 : _GEN_2012; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2014 = 8'hde == io_in_3 ? 8'h21 : _GEN_2013; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2015 = 8'hdf == io_in_3 ? 8'h2c : _GEN_2014; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2016 = 8'he0 == io_in_3 ? 8'hc : _GEN_2015; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2017 = 8'he1 == io_in_3 ? 8'h1 : _GEN_2016; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2018 = 8'he2 == io_in_3 ? 8'h16 : _GEN_2017; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2019 = 8'he3 == io_in_3 ? 8'h1b : _GEN_2018; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2020 = 8'he4 == io_in_3 ? 8'h38 : _GEN_2019; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2021 = 8'he5 == io_in_3 ? 8'h35 : _GEN_2020; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2022 = 8'he6 == io_in_3 ? 8'h22 : _GEN_2021; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2023 = 8'he7 == io_in_3 ? 8'h2f : _GEN_2022; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2024 = 8'he8 == io_in_3 ? 8'h64 : _GEN_2023; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2025 = 8'he9 == io_in_3 ? 8'h69 : _GEN_2024; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2026 = 8'hea == io_in_3 ? 8'h7e : _GEN_2025; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2027 = 8'heb == io_in_3 ? 8'h73 : _GEN_2026; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2028 = 8'hec == io_in_3 ? 8'h50 : _GEN_2027; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2029 = 8'hed == io_in_3 ? 8'h5d : _GEN_2028; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2030 = 8'hee == io_in_3 ? 8'h4a : _GEN_2029; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2031 = 8'hef == io_in_3 ? 8'h47 : _GEN_2030; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2032 = 8'hf0 == io_in_3 ? 8'hdc : _GEN_2031; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2033 = 8'hf1 == io_in_3 ? 8'hd1 : _GEN_2032; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2034 = 8'hf2 == io_in_3 ? 8'hc6 : _GEN_2033; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2035 = 8'hf3 == io_in_3 ? 8'hcb : _GEN_2034; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2036 = 8'hf4 == io_in_3 ? 8'he8 : _GEN_2035; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2037 = 8'hf5 == io_in_3 ? 8'he5 : _GEN_2036; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2038 = 8'hf6 == io_in_3 ? 8'hf2 : _GEN_2037; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2039 = 8'hf7 == io_in_3 ? 8'hff : _GEN_2038; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2040 = 8'hf8 == io_in_3 ? 8'hb4 : _GEN_2039; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2041 = 8'hf9 == io_in_3 ? 8'hb9 : _GEN_2040; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2042 = 8'hfa == io_in_3 ? 8'hae : _GEN_2041; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2043 = 8'hfb == io_in_3 ? 8'ha3 : _GEN_2042; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2044 = 8'hfc == io_in_3 ? 8'h80 : _GEN_2043; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2045 = 8'hfd == io_in_3 ? 8'h8d : _GEN_2044; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2046 = 8'hfe == io_in_3 ? 8'h9a : _GEN_2045; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2047 = 8'hff == io_in_3 ? 8'h97 : _GEN_2046; // @[AES_PipelinedElasticBuffer.scala 592:67 AES_PipelinedElasticBuffer.scala 592:67]
  wire [7:0] _GEN_2049 = 8'h1 == io_in_0 ? 8'hd : 8'h0; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2050 = 8'h2 == io_in_0 ? 8'h1a : _GEN_2049; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2051 = 8'h3 == io_in_0 ? 8'h17 : _GEN_2050; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2052 = 8'h4 == io_in_0 ? 8'h34 : _GEN_2051; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2053 = 8'h5 == io_in_0 ? 8'h39 : _GEN_2052; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2054 = 8'h6 == io_in_0 ? 8'h2e : _GEN_2053; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2055 = 8'h7 == io_in_0 ? 8'h23 : _GEN_2054; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2056 = 8'h8 == io_in_0 ? 8'h68 : _GEN_2055; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2057 = 8'h9 == io_in_0 ? 8'h65 : _GEN_2056; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2058 = 8'ha == io_in_0 ? 8'h72 : _GEN_2057; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2059 = 8'hb == io_in_0 ? 8'h7f : _GEN_2058; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2060 = 8'hc == io_in_0 ? 8'h5c : _GEN_2059; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2061 = 8'hd == io_in_0 ? 8'h51 : _GEN_2060; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2062 = 8'he == io_in_0 ? 8'h46 : _GEN_2061; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2063 = 8'hf == io_in_0 ? 8'h4b : _GEN_2062; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2064 = 8'h10 == io_in_0 ? 8'hd0 : _GEN_2063; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2065 = 8'h11 == io_in_0 ? 8'hdd : _GEN_2064; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2066 = 8'h12 == io_in_0 ? 8'hca : _GEN_2065; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2067 = 8'h13 == io_in_0 ? 8'hc7 : _GEN_2066; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2068 = 8'h14 == io_in_0 ? 8'he4 : _GEN_2067; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2069 = 8'h15 == io_in_0 ? 8'he9 : _GEN_2068; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2070 = 8'h16 == io_in_0 ? 8'hfe : _GEN_2069; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2071 = 8'h17 == io_in_0 ? 8'hf3 : _GEN_2070; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2072 = 8'h18 == io_in_0 ? 8'hb8 : _GEN_2071; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2073 = 8'h19 == io_in_0 ? 8'hb5 : _GEN_2072; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2074 = 8'h1a == io_in_0 ? 8'ha2 : _GEN_2073; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2075 = 8'h1b == io_in_0 ? 8'haf : _GEN_2074; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2076 = 8'h1c == io_in_0 ? 8'h8c : _GEN_2075; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2077 = 8'h1d == io_in_0 ? 8'h81 : _GEN_2076; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2078 = 8'h1e == io_in_0 ? 8'h96 : _GEN_2077; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2079 = 8'h1f == io_in_0 ? 8'h9b : _GEN_2078; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2080 = 8'h20 == io_in_0 ? 8'hbb : _GEN_2079; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2081 = 8'h21 == io_in_0 ? 8'hb6 : _GEN_2080; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2082 = 8'h22 == io_in_0 ? 8'ha1 : _GEN_2081; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2083 = 8'h23 == io_in_0 ? 8'hac : _GEN_2082; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2084 = 8'h24 == io_in_0 ? 8'h8f : _GEN_2083; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2085 = 8'h25 == io_in_0 ? 8'h82 : _GEN_2084; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2086 = 8'h26 == io_in_0 ? 8'h95 : _GEN_2085; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2087 = 8'h27 == io_in_0 ? 8'h98 : _GEN_2086; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2088 = 8'h28 == io_in_0 ? 8'hd3 : _GEN_2087; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2089 = 8'h29 == io_in_0 ? 8'hde : _GEN_2088; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2090 = 8'h2a == io_in_0 ? 8'hc9 : _GEN_2089; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2091 = 8'h2b == io_in_0 ? 8'hc4 : _GEN_2090; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2092 = 8'h2c == io_in_0 ? 8'he7 : _GEN_2091; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2093 = 8'h2d == io_in_0 ? 8'hea : _GEN_2092; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2094 = 8'h2e == io_in_0 ? 8'hfd : _GEN_2093; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2095 = 8'h2f == io_in_0 ? 8'hf0 : _GEN_2094; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2096 = 8'h30 == io_in_0 ? 8'h6b : _GEN_2095; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2097 = 8'h31 == io_in_0 ? 8'h66 : _GEN_2096; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2098 = 8'h32 == io_in_0 ? 8'h71 : _GEN_2097; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2099 = 8'h33 == io_in_0 ? 8'h7c : _GEN_2098; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2100 = 8'h34 == io_in_0 ? 8'h5f : _GEN_2099; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2101 = 8'h35 == io_in_0 ? 8'h52 : _GEN_2100; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2102 = 8'h36 == io_in_0 ? 8'h45 : _GEN_2101; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2103 = 8'h37 == io_in_0 ? 8'h48 : _GEN_2102; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2104 = 8'h38 == io_in_0 ? 8'h3 : _GEN_2103; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2105 = 8'h39 == io_in_0 ? 8'he : _GEN_2104; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2106 = 8'h3a == io_in_0 ? 8'h19 : _GEN_2105; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2107 = 8'h3b == io_in_0 ? 8'h14 : _GEN_2106; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2108 = 8'h3c == io_in_0 ? 8'h37 : _GEN_2107; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2109 = 8'h3d == io_in_0 ? 8'h3a : _GEN_2108; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2110 = 8'h3e == io_in_0 ? 8'h2d : _GEN_2109; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2111 = 8'h3f == io_in_0 ? 8'h20 : _GEN_2110; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2112 = 8'h40 == io_in_0 ? 8'h6d : _GEN_2111; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2113 = 8'h41 == io_in_0 ? 8'h60 : _GEN_2112; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2114 = 8'h42 == io_in_0 ? 8'h77 : _GEN_2113; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2115 = 8'h43 == io_in_0 ? 8'h7a : _GEN_2114; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2116 = 8'h44 == io_in_0 ? 8'h59 : _GEN_2115; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2117 = 8'h45 == io_in_0 ? 8'h54 : _GEN_2116; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2118 = 8'h46 == io_in_0 ? 8'h43 : _GEN_2117; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2119 = 8'h47 == io_in_0 ? 8'h4e : _GEN_2118; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2120 = 8'h48 == io_in_0 ? 8'h5 : _GEN_2119; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2121 = 8'h49 == io_in_0 ? 8'h8 : _GEN_2120; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2122 = 8'h4a == io_in_0 ? 8'h1f : _GEN_2121; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2123 = 8'h4b == io_in_0 ? 8'h12 : _GEN_2122; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2124 = 8'h4c == io_in_0 ? 8'h31 : _GEN_2123; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2125 = 8'h4d == io_in_0 ? 8'h3c : _GEN_2124; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2126 = 8'h4e == io_in_0 ? 8'h2b : _GEN_2125; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2127 = 8'h4f == io_in_0 ? 8'h26 : _GEN_2126; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2128 = 8'h50 == io_in_0 ? 8'hbd : _GEN_2127; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2129 = 8'h51 == io_in_0 ? 8'hb0 : _GEN_2128; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2130 = 8'h52 == io_in_0 ? 8'ha7 : _GEN_2129; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2131 = 8'h53 == io_in_0 ? 8'haa : _GEN_2130; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2132 = 8'h54 == io_in_0 ? 8'h89 : _GEN_2131; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2133 = 8'h55 == io_in_0 ? 8'h84 : _GEN_2132; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2134 = 8'h56 == io_in_0 ? 8'h93 : _GEN_2133; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2135 = 8'h57 == io_in_0 ? 8'h9e : _GEN_2134; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2136 = 8'h58 == io_in_0 ? 8'hd5 : _GEN_2135; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2137 = 8'h59 == io_in_0 ? 8'hd8 : _GEN_2136; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2138 = 8'h5a == io_in_0 ? 8'hcf : _GEN_2137; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2139 = 8'h5b == io_in_0 ? 8'hc2 : _GEN_2138; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2140 = 8'h5c == io_in_0 ? 8'he1 : _GEN_2139; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2141 = 8'h5d == io_in_0 ? 8'hec : _GEN_2140; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2142 = 8'h5e == io_in_0 ? 8'hfb : _GEN_2141; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2143 = 8'h5f == io_in_0 ? 8'hf6 : _GEN_2142; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2144 = 8'h60 == io_in_0 ? 8'hd6 : _GEN_2143; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2145 = 8'h61 == io_in_0 ? 8'hdb : _GEN_2144; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2146 = 8'h62 == io_in_0 ? 8'hcc : _GEN_2145; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2147 = 8'h63 == io_in_0 ? 8'hc1 : _GEN_2146; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2148 = 8'h64 == io_in_0 ? 8'he2 : _GEN_2147; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2149 = 8'h65 == io_in_0 ? 8'hef : _GEN_2148; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2150 = 8'h66 == io_in_0 ? 8'hf8 : _GEN_2149; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2151 = 8'h67 == io_in_0 ? 8'hf5 : _GEN_2150; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2152 = 8'h68 == io_in_0 ? 8'hbe : _GEN_2151; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2153 = 8'h69 == io_in_0 ? 8'hb3 : _GEN_2152; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2154 = 8'h6a == io_in_0 ? 8'ha4 : _GEN_2153; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2155 = 8'h6b == io_in_0 ? 8'ha9 : _GEN_2154; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2156 = 8'h6c == io_in_0 ? 8'h8a : _GEN_2155; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2157 = 8'h6d == io_in_0 ? 8'h87 : _GEN_2156; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2158 = 8'h6e == io_in_0 ? 8'h90 : _GEN_2157; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2159 = 8'h6f == io_in_0 ? 8'h9d : _GEN_2158; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2160 = 8'h70 == io_in_0 ? 8'h6 : _GEN_2159; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2161 = 8'h71 == io_in_0 ? 8'hb : _GEN_2160; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2162 = 8'h72 == io_in_0 ? 8'h1c : _GEN_2161; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2163 = 8'h73 == io_in_0 ? 8'h11 : _GEN_2162; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2164 = 8'h74 == io_in_0 ? 8'h32 : _GEN_2163; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2165 = 8'h75 == io_in_0 ? 8'h3f : _GEN_2164; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2166 = 8'h76 == io_in_0 ? 8'h28 : _GEN_2165; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2167 = 8'h77 == io_in_0 ? 8'h25 : _GEN_2166; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2168 = 8'h78 == io_in_0 ? 8'h6e : _GEN_2167; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2169 = 8'h79 == io_in_0 ? 8'h63 : _GEN_2168; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2170 = 8'h7a == io_in_0 ? 8'h74 : _GEN_2169; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2171 = 8'h7b == io_in_0 ? 8'h79 : _GEN_2170; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2172 = 8'h7c == io_in_0 ? 8'h5a : _GEN_2171; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2173 = 8'h7d == io_in_0 ? 8'h57 : _GEN_2172; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2174 = 8'h7e == io_in_0 ? 8'h40 : _GEN_2173; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2175 = 8'h7f == io_in_0 ? 8'h4d : _GEN_2174; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2176 = 8'h80 == io_in_0 ? 8'hda : _GEN_2175; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2177 = 8'h81 == io_in_0 ? 8'hd7 : _GEN_2176; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2178 = 8'h82 == io_in_0 ? 8'hc0 : _GEN_2177; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2179 = 8'h83 == io_in_0 ? 8'hcd : _GEN_2178; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2180 = 8'h84 == io_in_0 ? 8'hee : _GEN_2179; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2181 = 8'h85 == io_in_0 ? 8'he3 : _GEN_2180; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2182 = 8'h86 == io_in_0 ? 8'hf4 : _GEN_2181; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2183 = 8'h87 == io_in_0 ? 8'hf9 : _GEN_2182; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2184 = 8'h88 == io_in_0 ? 8'hb2 : _GEN_2183; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2185 = 8'h89 == io_in_0 ? 8'hbf : _GEN_2184; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2186 = 8'h8a == io_in_0 ? 8'ha8 : _GEN_2185; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2187 = 8'h8b == io_in_0 ? 8'ha5 : _GEN_2186; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2188 = 8'h8c == io_in_0 ? 8'h86 : _GEN_2187; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2189 = 8'h8d == io_in_0 ? 8'h8b : _GEN_2188; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2190 = 8'h8e == io_in_0 ? 8'h9c : _GEN_2189; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2191 = 8'h8f == io_in_0 ? 8'h91 : _GEN_2190; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2192 = 8'h90 == io_in_0 ? 8'ha : _GEN_2191; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2193 = 8'h91 == io_in_0 ? 8'h7 : _GEN_2192; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2194 = 8'h92 == io_in_0 ? 8'h10 : _GEN_2193; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2195 = 8'h93 == io_in_0 ? 8'h1d : _GEN_2194; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2196 = 8'h94 == io_in_0 ? 8'h3e : _GEN_2195; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2197 = 8'h95 == io_in_0 ? 8'h33 : _GEN_2196; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2198 = 8'h96 == io_in_0 ? 8'h24 : _GEN_2197; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2199 = 8'h97 == io_in_0 ? 8'h29 : _GEN_2198; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2200 = 8'h98 == io_in_0 ? 8'h62 : _GEN_2199; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2201 = 8'h99 == io_in_0 ? 8'h6f : _GEN_2200; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2202 = 8'h9a == io_in_0 ? 8'h78 : _GEN_2201; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2203 = 8'h9b == io_in_0 ? 8'h75 : _GEN_2202; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2204 = 8'h9c == io_in_0 ? 8'h56 : _GEN_2203; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2205 = 8'h9d == io_in_0 ? 8'h5b : _GEN_2204; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2206 = 8'h9e == io_in_0 ? 8'h4c : _GEN_2205; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2207 = 8'h9f == io_in_0 ? 8'h41 : _GEN_2206; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2208 = 8'ha0 == io_in_0 ? 8'h61 : _GEN_2207; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2209 = 8'ha1 == io_in_0 ? 8'h6c : _GEN_2208; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2210 = 8'ha2 == io_in_0 ? 8'h7b : _GEN_2209; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2211 = 8'ha3 == io_in_0 ? 8'h76 : _GEN_2210; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2212 = 8'ha4 == io_in_0 ? 8'h55 : _GEN_2211; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2213 = 8'ha5 == io_in_0 ? 8'h58 : _GEN_2212; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2214 = 8'ha6 == io_in_0 ? 8'h4f : _GEN_2213; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2215 = 8'ha7 == io_in_0 ? 8'h42 : _GEN_2214; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2216 = 8'ha8 == io_in_0 ? 8'h9 : _GEN_2215; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2217 = 8'ha9 == io_in_0 ? 8'h4 : _GEN_2216; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2218 = 8'haa == io_in_0 ? 8'h13 : _GEN_2217; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2219 = 8'hab == io_in_0 ? 8'h1e : _GEN_2218; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2220 = 8'hac == io_in_0 ? 8'h3d : _GEN_2219; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2221 = 8'had == io_in_0 ? 8'h30 : _GEN_2220; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2222 = 8'hae == io_in_0 ? 8'h27 : _GEN_2221; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2223 = 8'haf == io_in_0 ? 8'h2a : _GEN_2222; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2224 = 8'hb0 == io_in_0 ? 8'hb1 : _GEN_2223; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2225 = 8'hb1 == io_in_0 ? 8'hbc : _GEN_2224; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2226 = 8'hb2 == io_in_0 ? 8'hab : _GEN_2225; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2227 = 8'hb3 == io_in_0 ? 8'ha6 : _GEN_2226; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2228 = 8'hb4 == io_in_0 ? 8'h85 : _GEN_2227; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2229 = 8'hb5 == io_in_0 ? 8'h88 : _GEN_2228; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2230 = 8'hb6 == io_in_0 ? 8'h9f : _GEN_2229; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2231 = 8'hb7 == io_in_0 ? 8'h92 : _GEN_2230; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2232 = 8'hb8 == io_in_0 ? 8'hd9 : _GEN_2231; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2233 = 8'hb9 == io_in_0 ? 8'hd4 : _GEN_2232; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2234 = 8'hba == io_in_0 ? 8'hc3 : _GEN_2233; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2235 = 8'hbb == io_in_0 ? 8'hce : _GEN_2234; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2236 = 8'hbc == io_in_0 ? 8'hed : _GEN_2235; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2237 = 8'hbd == io_in_0 ? 8'he0 : _GEN_2236; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2238 = 8'hbe == io_in_0 ? 8'hf7 : _GEN_2237; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2239 = 8'hbf == io_in_0 ? 8'hfa : _GEN_2238; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2240 = 8'hc0 == io_in_0 ? 8'hb7 : _GEN_2239; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2241 = 8'hc1 == io_in_0 ? 8'hba : _GEN_2240; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2242 = 8'hc2 == io_in_0 ? 8'had : _GEN_2241; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2243 = 8'hc3 == io_in_0 ? 8'ha0 : _GEN_2242; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2244 = 8'hc4 == io_in_0 ? 8'h83 : _GEN_2243; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2245 = 8'hc5 == io_in_0 ? 8'h8e : _GEN_2244; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2246 = 8'hc6 == io_in_0 ? 8'h99 : _GEN_2245; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2247 = 8'hc7 == io_in_0 ? 8'h94 : _GEN_2246; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2248 = 8'hc8 == io_in_0 ? 8'hdf : _GEN_2247; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2249 = 8'hc9 == io_in_0 ? 8'hd2 : _GEN_2248; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2250 = 8'hca == io_in_0 ? 8'hc5 : _GEN_2249; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2251 = 8'hcb == io_in_0 ? 8'hc8 : _GEN_2250; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2252 = 8'hcc == io_in_0 ? 8'heb : _GEN_2251; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2253 = 8'hcd == io_in_0 ? 8'he6 : _GEN_2252; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2254 = 8'hce == io_in_0 ? 8'hf1 : _GEN_2253; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2255 = 8'hcf == io_in_0 ? 8'hfc : _GEN_2254; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2256 = 8'hd0 == io_in_0 ? 8'h67 : _GEN_2255; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2257 = 8'hd1 == io_in_0 ? 8'h6a : _GEN_2256; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2258 = 8'hd2 == io_in_0 ? 8'h7d : _GEN_2257; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2259 = 8'hd3 == io_in_0 ? 8'h70 : _GEN_2258; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2260 = 8'hd4 == io_in_0 ? 8'h53 : _GEN_2259; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2261 = 8'hd5 == io_in_0 ? 8'h5e : _GEN_2260; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2262 = 8'hd6 == io_in_0 ? 8'h49 : _GEN_2261; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2263 = 8'hd7 == io_in_0 ? 8'h44 : _GEN_2262; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2264 = 8'hd8 == io_in_0 ? 8'hf : _GEN_2263; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2265 = 8'hd9 == io_in_0 ? 8'h2 : _GEN_2264; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2266 = 8'hda == io_in_0 ? 8'h15 : _GEN_2265; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2267 = 8'hdb == io_in_0 ? 8'h18 : _GEN_2266; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2268 = 8'hdc == io_in_0 ? 8'h3b : _GEN_2267; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2269 = 8'hdd == io_in_0 ? 8'h36 : _GEN_2268; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2270 = 8'hde == io_in_0 ? 8'h21 : _GEN_2269; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2271 = 8'hdf == io_in_0 ? 8'h2c : _GEN_2270; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2272 = 8'he0 == io_in_0 ? 8'hc : _GEN_2271; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2273 = 8'he1 == io_in_0 ? 8'h1 : _GEN_2272; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2274 = 8'he2 == io_in_0 ? 8'h16 : _GEN_2273; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2275 = 8'he3 == io_in_0 ? 8'h1b : _GEN_2274; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2276 = 8'he4 == io_in_0 ? 8'h38 : _GEN_2275; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2277 = 8'he5 == io_in_0 ? 8'h35 : _GEN_2276; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2278 = 8'he6 == io_in_0 ? 8'h22 : _GEN_2277; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2279 = 8'he7 == io_in_0 ? 8'h2f : _GEN_2278; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2280 = 8'he8 == io_in_0 ? 8'h64 : _GEN_2279; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2281 = 8'he9 == io_in_0 ? 8'h69 : _GEN_2280; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2282 = 8'hea == io_in_0 ? 8'h7e : _GEN_2281; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2283 = 8'heb == io_in_0 ? 8'h73 : _GEN_2282; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2284 = 8'hec == io_in_0 ? 8'h50 : _GEN_2283; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2285 = 8'hed == io_in_0 ? 8'h5d : _GEN_2284; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2286 = 8'hee == io_in_0 ? 8'h4a : _GEN_2285; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2287 = 8'hef == io_in_0 ? 8'h47 : _GEN_2286; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2288 = 8'hf0 == io_in_0 ? 8'hdc : _GEN_2287; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2289 = 8'hf1 == io_in_0 ? 8'hd1 : _GEN_2288; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2290 = 8'hf2 == io_in_0 ? 8'hc6 : _GEN_2289; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2291 = 8'hf3 == io_in_0 ? 8'hcb : _GEN_2290; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2292 = 8'hf4 == io_in_0 ? 8'he8 : _GEN_2291; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2293 = 8'hf5 == io_in_0 ? 8'he5 : _GEN_2292; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2294 = 8'hf6 == io_in_0 ? 8'hf2 : _GEN_2293; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2295 = 8'hf7 == io_in_0 ? 8'hff : _GEN_2294; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2296 = 8'hf8 == io_in_0 ? 8'hb4 : _GEN_2295; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2297 = 8'hf9 == io_in_0 ? 8'hb9 : _GEN_2296; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2298 = 8'hfa == io_in_0 ? 8'hae : _GEN_2297; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2299 = 8'hfb == io_in_0 ? 8'ha3 : _GEN_2298; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2300 = 8'hfc == io_in_0 ? 8'h80 : _GEN_2299; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2301 = 8'hfd == io_in_0 ? 8'h8d : _GEN_2300; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2302 = 8'hfe == io_in_0 ? 8'h9a : _GEN_2301; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2303 = 8'hff == io_in_0 ? 8'h97 : _GEN_2302; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2305 = 8'h1 == io_in_1 ? 8'h9 : 8'h0; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2306 = 8'h2 == io_in_1 ? 8'h12 : _GEN_2305; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2307 = 8'h3 == io_in_1 ? 8'h1b : _GEN_2306; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2308 = 8'h4 == io_in_1 ? 8'h24 : _GEN_2307; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2309 = 8'h5 == io_in_1 ? 8'h2d : _GEN_2308; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2310 = 8'h6 == io_in_1 ? 8'h36 : _GEN_2309; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2311 = 8'h7 == io_in_1 ? 8'h3f : _GEN_2310; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2312 = 8'h8 == io_in_1 ? 8'h48 : _GEN_2311; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2313 = 8'h9 == io_in_1 ? 8'h41 : _GEN_2312; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2314 = 8'ha == io_in_1 ? 8'h5a : _GEN_2313; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2315 = 8'hb == io_in_1 ? 8'h53 : _GEN_2314; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2316 = 8'hc == io_in_1 ? 8'h6c : _GEN_2315; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2317 = 8'hd == io_in_1 ? 8'h65 : _GEN_2316; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2318 = 8'he == io_in_1 ? 8'h7e : _GEN_2317; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2319 = 8'hf == io_in_1 ? 8'h77 : _GEN_2318; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2320 = 8'h10 == io_in_1 ? 8'h90 : _GEN_2319; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2321 = 8'h11 == io_in_1 ? 8'h99 : _GEN_2320; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2322 = 8'h12 == io_in_1 ? 8'h82 : _GEN_2321; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2323 = 8'h13 == io_in_1 ? 8'h8b : _GEN_2322; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2324 = 8'h14 == io_in_1 ? 8'hb4 : _GEN_2323; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2325 = 8'h15 == io_in_1 ? 8'hbd : _GEN_2324; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2326 = 8'h16 == io_in_1 ? 8'ha6 : _GEN_2325; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2327 = 8'h17 == io_in_1 ? 8'haf : _GEN_2326; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2328 = 8'h18 == io_in_1 ? 8'hd8 : _GEN_2327; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2329 = 8'h19 == io_in_1 ? 8'hd1 : _GEN_2328; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2330 = 8'h1a == io_in_1 ? 8'hca : _GEN_2329; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2331 = 8'h1b == io_in_1 ? 8'hc3 : _GEN_2330; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2332 = 8'h1c == io_in_1 ? 8'hfc : _GEN_2331; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2333 = 8'h1d == io_in_1 ? 8'hf5 : _GEN_2332; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2334 = 8'h1e == io_in_1 ? 8'hee : _GEN_2333; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2335 = 8'h1f == io_in_1 ? 8'he7 : _GEN_2334; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2336 = 8'h20 == io_in_1 ? 8'h3b : _GEN_2335; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2337 = 8'h21 == io_in_1 ? 8'h32 : _GEN_2336; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2338 = 8'h22 == io_in_1 ? 8'h29 : _GEN_2337; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2339 = 8'h23 == io_in_1 ? 8'h20 : _GEN_2338; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2340 = 8'h24 == io_in_1 ? 8'h1f : _GEN_2339; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2341 = 8'h25 == io_in_1 ? 8'h16 : _GEN_2340; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2342 = 8'h26 == io_in_1 ? 8'hd : _GEN_2341; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2343 = 8'h27 == io_in_1 ? 8'h4 : _GEN_2342; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2344 = 8'h28 == io_in_1 ? 8'h73 : _GEN_2343; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2345 = 8'h29 == io_in_1 ? 8'h7a : _GEN_2344; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2346 = 8'h2a == io_in_1 ? 8'h61 : _GEN_2345; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2347 = 8'h2b == io_in_1 ? 8'h68 : _GEN_2346; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2348 = 8'h2c == io_in_1 ? 8'h57 : _GEN_2347; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2349 = 8'h2d == io_in_1 ? 8'h5e : _GEN_2348; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2350 = 8'h2e == io_in_1 ? 8'h45 : _GEN_2349; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2351 = 8'h2f == io_in_1 ? 8'h4c : _GEN_2350; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2352 = 8'h30 == io_in_1 ? 8'hab : _GEN_2351; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2353 = 8'h31 == io_in_1 ? 8'ha2 : _GEN_2352; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2354 = 8'h32 == io_in_1 ? 8'hb9 : _GEN_2353; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2355 = 8'h33 == io_in_1 ? 8'hb0 : _GEN_2354; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2356 = 8'h34 == io_in_1 ? 8'h8f : _GEN_2355; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2357 = 8'h35 == io_in_1 ? 8'h86 : _GEN_2356; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2358 = 8'h36 == io_in_1 ? 8'h9d : _GEN_2357; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2359 = 8'h37 == io_in_1 ? 8'h94 : _GEN_2358; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2360 = 8'h38 == io_in_1 ? 8'he3 : _GEN_2359; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2361 = 8'h39 == io_in_1 ? 8'hea : _GEN_2360; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2362 = 8'h3a == io_in_1 ? 8'hf1 : _GEN_2361; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2363 = 8'h3b == io_in_1 ? 8'hf8 : _GEN_2362; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2364 = 8'h3c == io_in_1 ? 8'hc7 : _GEN_2363; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2365 = 8'h3d == io_in_1 ? 8'hce : _GEN_2364; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2366 = 8'h3e == io_in_1 ? 8'hd5 : _GEN_2365; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2367 = 8'h3f == io_in_1 ? 8'hdc : _GEN_2366; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2368 = 8'h40 == io_in_1 ? 8'h76 : _GEN_2367; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2369 = 8'h41 == io_in_1 ? 8'h7f : _GEN_2368; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2370 = 8'h42 == io_in_1 ? 8'h64 : _GEN_2369; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2371 = 8'h43 == io_in_1 ? 8'h6d : _GEN_2370; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2372 = 8'h44 == io_in_1 ? 8'h52 : _GEN_2371; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2373 = 8'h45 == io_in_1 ? 8'h5b : _GEN_2372; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2374 = 8'h46 == io_in_1 ? 8'h40 : _GEN_2373; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2375 = 8'h47 == io_in_1 ? 8'h49 : _GEN_2374; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2376 = 8'h48 == io_in_1 ? 8'h3e : _GEN_2375; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2377 = 8'h49 == io_in_1 ? 8'h37 : _GEN_2376; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2378 = 8'h4a == io_in_1 ? 8'h2c : _GEN_2377; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2379 = 8'h4b == io_in_1 ? 8'h25 : _GEN_2378; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2380 = 8'h4c == io_in_1 ? 8'h1a : _GEN_2379; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2381 = 8'h4d == io_in_1 ? 8'h13 : _GEN_2380; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2382 = 8'h4e == io_in_1 ? 8'h8 : _GEN_2381; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2383 = 8'h4f == io_in_1 ? 8'h1 : _GEN_2382; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2384 = 8'h50 == io_in_1 ? 8'he6 : _GEN_2383; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2385 = 8'h51 == io_in_1 ? 8'hef : _GEN_2384; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2386 = 8'h52 == io_in_1 ? 8'hf4 : _GEN_2385; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2387 = 8'h53 == io_in_1 ? 8'hfd : _GEN_2386; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2388 = 8'h54 == io_in_1 ? 8'hc2 : _GEN_2387; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2389 = 8'h55 == io_in_1 ? 8'hcb : _GEN_2388; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2390 = 8'h56 == io_in_1 ? 8'hd0 : _GEN_2389; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2391 = 8'h57 == io_in_1 ? 8'hd9 : _GEN_2390; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2392 = 8'h58 == io_in_1 ? 8'hae : _GEN_2391; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2393 = 8'h59 == io_in_1 ? 8'ha7 : _GEN_2392; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2394 = 8'h5a == io_in_1 ? 8'hbc : _GEN_2393; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2395 = 8'h5b == io_in_1 ? 8'hb5 : _GEN_2394; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2396 = 8'h5c == io_in_1 ? 8'h8a : _GEN_2395; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2397 = 8'h5d == io_in_1 ? 8'h83 : _GEN_2396; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2398 = 8'h5e == io_in_1 ? 8'h98 : _GEN_2397; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2399 = 8'h5f == io_in_1 ? 8'h91 : _GEN_2398; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2400 = 8'h60 == io_in_1 ? 8'h4d : _GEN_2399; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2401 = 8'h61 == io_in_1 ? 8'h44 : _GEN_2400; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2402 = 8'h62 == io_in_1 ? 8'h5f : _GEN_2401; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2403 = 8'h63 == io_in_1 ? 8'h56 : _GEN_2402; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2404 = 8'h64 == io_in_1 ? 8'h69 : _GEN_2403; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2405 = 8'h65 == io_in_1 ? 8'h60 : _GEN_2404; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2406 = 8'h66 == io_in_1 ? 8'h7b : _GEN_2405; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2407 = 8'h67 == io_in_1 ? 8'h72 : _GEN_2406; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2408 = 8'h68 == io_in_1 ? 8'h5 : _GEN_2407; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2409 = 8'h69 == io_in_1 ? 8'hc : _GEN_2408; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2410 = 8'h6a == io_in_1 ? 8'h17 : _GEN_2409; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2411 = 8'h6b == io_in_1 ? 8'h1e : _GEN_2410; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2412 = 8'h6c == io_in_1 ? 8'h21 : _GEN_2411; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2413 = 8'h6d == io_in_1 ? 8'h28 : _GEN_2412; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2414 = 8'h6e == io_in_1 ? 8'h33 : _GEN_2413; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2415 = 8'h6f == io_in_1 ? 8'h3a : _GEN_2414; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2416 = 8'h70 == io_in_1 ? 8'hdd : _GEN_2415; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2417 = 8'h71 == io_in_1 ? 8'hd4 : _GEN_2416; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2418 = 8'h72 == io_in_1 ? 8'hcf : _GEN_2417; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2419 = 8'h73 == io_in_1 ? 8'hc6 : _GEN_2418; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2420 = 8'h74 == io_in_1 ? 8'hf9 : _GEN_2419; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2421 = 8'h75 == io_in_1 ? 8'hf0 : _GEN_2420; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2422 = 8'h76 == io_in_1 ? 8'heb : _GEN_2421; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2423 = 8'h77 == io_in_1 ? 8'he2 : _GEN_2422; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2424 = 8'h78 == io_in_1 ? 8'h95 : _GEN_2423; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2425 = 8'h79 == io_in_1 ? 8'h9c : _GEN_2424; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2426 = 8'h7a == io_in_1 ? 8'h87 : _GEN_2425; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2427 = 8'h7b == io_in_1 ? 8'h8e : _GEN_2426; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2428 = 8'h7c == io_in_1 ? 8'hb1 : _GEN_2427; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2429 = 8'h7d == io_in_1 ? 8'hb8 : _GEN_2428; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2430 = 8'h7e == io_in_1 ? 8'ha3 : _GEN_2429; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2431 = 8'h7f == io_in_1 ? 8'haa : _GEN_2430; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2432 = 8'h80 == io_in_1 ? 8'hec : _GEN_2431; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2433 = 8'h81 == io_in_1 ? 8'he5 : _GEN_2432; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2434 = 8'h82 == io_in_1 ? 8'hfe : _GEN_2433; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2435 = 8'h83 == io_in_1 ? 8'hf7 : _GEN_2434; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2436 = 8'h84 == io_in_1 ? 8'hc8 : _GEN_2435; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2437 = 8'h85 == io_in_1 ? 8'hc1 : _GEN_2436; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2438 = 8'h86 == io_in_1 ? 8'hda : _GEN_2437; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2439 = 8'h87 == io_in_1 ? 8'hd3 : _GEN_2438; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2440 = 8'h88 == io_in_1 ? 8'ha4 : _GEN_2439; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2441 = 8'h89 == io_in_1 ? 8'had : _GEN_2440; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2442 = 8'h8a == io_in_1 ? 8'hb6 : _GEN_2441; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2443 = 8'h8b == io_in_1 ? 8'hbf : _GEN_2442; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2444 = 8'h8c == io_in_1 ? 8'h80 : _GEN_2443; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2445 = 8'h8d == io_in_1 ? 8'h89 : _GEN_2444; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2446 = 8'h8e == io_in_1 ? 8'h92 : _GEN_2445; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2447 = 8'h8f == io_in_1 ? 8'h9b : _GEN_2446; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2448 = 8'h90 == io_in_1 ? 8'h7c : _GEN_2447; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2449 = 8'h91 == io_in_1 ? 8'h75 : _GEN_2448; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2450 = 8'h92 == io_in_1 ? 8'h6e : _GEN_2449; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2451 = 8'h93 == io_in_1 ? 8'h67 : _GEN_2450; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2452 = 8'h94 == io_in_1 ? 8'h58 : _GEN_2451; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2453 = 8'h95 == io_in_1 ? 8'h51 : _GEN_2452; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2454 = 8'h96 == io_in_1 ? 8'h4a : _GEN_2453; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2455 = 8'h97 == io_in_1 ? 8'h43 : _GEN_2454; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2456 = 8'h98 == io_in_1 ? 8'h34 : _GEN_2455; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2457 = 8'h99 == io_in_1 ? 8'h3d : _GEN_2456; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2458 = 8'h9a == io_in_1 ? 8'h26 : _GEN_2457; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2459 = 8'h9b == io_in_1 ? 8'h2f : _GEN_2458; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2460 = 8'h9c == io_in_1 ? 8'h10 : _GEN_2459; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2461 = 8'h9d == io_in_1 ? 8'h19 : _GEN_2460; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2462 = 8'h9e == io_in_1 ? 8'h2 : _GEN_2461; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2463 = 8'h9f == io_in_1 ? 8'hb : _GEN_2462; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2464 = 8'ha0 == io_in_1 ? 8'hd7 : _GEN_2463; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2465 = 8'ha1 == io_in_1 ? 8'hde : _GEN_2464; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2466 = 8'ha2 == io_in_1 ? 8'hc5 : _GEN_2465; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2467 = 8'ha3 == io_in_1 ? 8'hcc : _GEN_2466; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2468 = 8'ha4 == io_in_1 ? 8'hf3 : _GEN_2467; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2469 = 8'ha5 == io_in_1 ? 8'hfa : _GEN_2468; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2470 = 8'ha6 == io_in_1 ? 8'he1 : _GEN_2469; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2471 = 8'ha7 == io_in_1 ? 8'he8 : _GEN_2470; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2472 = 8'ha8 == io_in_1 ? 8'h9f : _GEN_2471; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2473 = 8'ha9 == io_in_1 ? 8'h96 : _GEN_2472; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2474 = 8'haa == io_in_1 ? 8'h8d : _GEN_2473; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2475 = 8'hab == io_in_1 ? 8'h84 : _GEN_2474; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2476 = 8'hac == io_in_1 ? 8'hbb : _GEN_2475; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2477 = 8'had == io_in_1 ? 8'hb2 : _GEN_2476; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2478 = 8'hae == io_in_1 ? 8'ha9 : _GEN_2477; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2479 = 8'haf == io_in_1 ? 8'ha0 : _GEN_2478; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2480 = 8'hb0 == io_in_1 ? 8'h47 : _GEN_2479; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2481 = 8'hb1 == io_in_1 ? 8'h4e : _GEN_2480; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2482 = 8'hb2 == io_in_1 ? 8'h55 : _GEN_2481; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2483 = 8'hb3 == io_in_1 ? 8'h5c : _GEN_2482; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2484 = 8'hb4 == io_in_1 ? 8'h63 : _GEN_2483; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2485 = 8'hb5 == io_in_1 ? 8'h6a : _GEN_2484; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2486 = 8'hb6 == io_in_1 ? 8'h71 : _GEN_2485; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2487 = 8'hb7 == io_in_1 ? 8'h78 : _GEN_2486; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2488 = 8'hb8 == io_in_1 ? 8'hf : _GEN_2487; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2489 = 8'hb9 == io_in_1 ? 8'h6 : _GEN_2488; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2490 = 8'hba == io_in_1 ? 8'h1d : _GEN_2489; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2491 = 8'hbb == io_in_1 ? 8'h14 : _GEN_2490; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2492 = 8'hbc == io_in_1 ? 8'h2b : _GEN_2491; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2493 = 8'hbd == io_in_1 ? 8'h22 : _GEN_2492; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2494 = 8'hbe == io_in_1 ? 8'h39 : _GEN_2493; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2495 = 8'hbf == io_in_1 ? 8'h30 : _GEN_2494; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2496 = 8'hc0 == io_in_1 ? 8'h9a : _GEN_2495; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2497 = 8'hc1 == io_in_1 ? 8'h93 : _GEN_2496; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2498 = 8'hc2 == io_in_1 ? 8'h88 : _GEN_2497; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2499 = 8'hc3 == io_in_1 ? 8'h81 : _GEN_2498; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2500 = 8'hc4 == io_in_1 ? 8'hbe : _GEN_2499; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2501 = 8'hc5 == io_in_1 ? 8'hb7 : _GEN_2500; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2502 = 8'hc6 == io_in_1 ? 8'hac : _GEN_2501; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2503 = 8'hc7 == io_in_1 ? 8'ha5 : _GEN_2502; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2504 = 8'hc8 == io_in_1 ? 8'hd2 : _GEN_2503; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2505 = 8'hc9 == io_in_1 ? 8'hdb : _GEN_2504; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2506 = 8'hca == io_in_1 ? 8'hc0 : _GEN_2505; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2507 = 8'hcb == io_in_1 ? 8'hc9 : _GEN_2506; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2508 = 8'hcc == io_in_1 ? 8'hf6 : _GEN_2507; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2509 = 8'hcd == io_in_1 ? 8'hff : _GEN_2508; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2510 = 8'hce == io_in_1 ? 8'he4 : _GEN_2509; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2511 = 8'hcf == io_in_1 ? 8'hed : _GEN_2510; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2512 = 8'hd0 == io_in_1 ? 8'ha : _GEN_2511; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2513 = 8'hd1 == io_in_1 ? 8'h3 : _GEN_2512; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2514 = 8'hd2 == io_in_1 ? 8'h18 : _GEN_2513; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2515 = 8'hd3 == io_in_1 ? 8'h11 : _GEN_2514; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2516 = 8'hd4 == io_in_1 ? 8'h2e : _GEN_2515; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2517 = 8'hd5 == io_in_1 ? 8'h27 : _GEN_2516; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2518 = 8'hd6 == io_in_1 ? 8'h3c : _GEN_2517; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2519 = 8'hd7 == io_in_1 ? 8'h35 : _GEN_2518; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2520 = 8'hd8 == io_in_1 ? 8'h42 : _GEN_2519; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2521 = 8'hd9 == io_in_1 ? 8'h4b : _GEN_2520; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2522 = 8'hda == io_in_1 ? 8'h50 : _GEN_2521; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2523 = 8'hdb == io_in_1 ? 8'h59 : _GEN_2522; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2524 = 8'hdc == io_in_1 ? 8'h66 : _GEN_2523; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2525 = 8'hdd == io_in_1 ? 8'h6f : _GEN_2524; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2526 = 8'hde == io_in_1 ? 8'h74 : _GEN_2525; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2527 = 8'hdf == io_in_1 ? 8'h7d : _GEN_2526; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2528 = 8'he0 == io_in_1 ? 8'ha1 : _GEN_2527; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2529 = 8'he1 == io_in_1 ? 8'ha8 : _GEN_2528; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2530 = 8'he2 == io_in_1 ? 8'hb3 : _GEN_2529; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2531 = 8'he3 == io_in_1 ? 8'hba : _GEN_2530; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2532 = 8'he4 == io_in_1 ? 8'h85 : _GEN_2531; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2533 = 8'he5 == io_in_1 ? 8'h8c : _GEN_2532; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2534 = 8'he6 == io_in_1 ? 8'h97 : _GEN_2533; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2535 = 8'he7 == io_in_1 ? 8'h9e : _GEN_2534; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2536 = 8'he8 == io_in_1 ? 8'he9 : _GEN_2535; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2537 = 8'he9 == io_in_1 ? 8'he0 : _GEN_2536; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2538 = 8'hea == io_in_1 ? 8'hfb : _GEN_2537; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2539 = 8'heb == io_in_1 ? 8'hf2 : _GEN_2538; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2540 = 8'hec == io_in_1 ? 8'hcd : _GEN_2539; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2541 = 8'hed == io_in_1 ? 8'hc4 : _GEN_2540; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2542 = 8'hee == io_in_1 ? 8'hdf : _GEN_2541; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2543 = 8'hef == io_in_1 ? 8'hd6 : _GEN_2542; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2544 = 8'hf0 == io_in_1 ? 8'h31 : _GEN_2543; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2545 = 8'hf1 == io_in_1 ? 8'h38 : _GEN_2544; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2546 = 8'hf2 == io_in_1 ? 8'h23 : _GEN_2545; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2547 = 8'hf3 == io_in_1 ? 8'h2a : _GEN_2546; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2548 = 8'hf4 == io_in_1 ? 8'h15 : _GEN_2547; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2549 = 8'hf5 == io_in_1 ? 8'h1c : _GEN_2548; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2550 = 8'hf6 == io_in_1 ? 8'h7 : _GEN_2549; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2551 = 8'hf7 == io_in_1 ? 8'he : _GEN_2550; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2552 = 8'hf8 == io_in_1 ? 8'h79 : _GEN_2551; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2553 = 8'hf9 == io_in_1 ? 8'h70 : _GEN_2552; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2554 = 8'hfa == io_in_1 ? 8'h6b : _GEN_2553; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2555 = 8'hfb == io_in_1 ? 8'h62 : _GEN_2554; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2556 = 8'hfc == io_in_1 ? 8'h5d : _GEN_2555; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2557 = 8'hfd == io_in_1 ? 8'h54 : _GEN_2556; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2558 = 8'hfe == io_in_1 ? 8'h4f : _GEN_2557; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2559 = 8'hff == io_in_1 ? 8'h46 : _GEN_2558; // @[AES_PipelinedElasticBuffer.scala 593:32 AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _T_6 = _GEN_2303 ^ _GEN_2559; // @[AES_PipelinedElasticBuffer.scala 593:32]
  wire [7:0] _GEN_2561 = 8'h1 == io_in_2 ? 8'he : 8'h0; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2562 = 8'h2 == io_in_2 ? 8'h1c : _GEN_2561; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2563 = 8'h3 == io_in_2 ? 8'h12 : _GEN_2562; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2564 = 8'h4 == io_in_2 ? 8'h38 : _GEN_2563; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2565 = 8'h5 == io_in_2 ? 8'h36 : _GEN_2564; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2566 = 8'h6 == io_in_2 ? 8'h24 : _GEN_2565; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2567 = 8'h7 == io_in_2 ? 8'h2a : _GEN_2566; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2568 = 8'h8 == io_in_2 ? 8'h70 : _GEN_2567; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2569 = 8'h9 == io_in_2 ? 8'h7e : _GEN_2568; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2570 = 8'ha == io_in_2 ? 8'h6c : _GEN_2569; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2571 = 8'hb == io_in_2 ? 8'h62 : _GEN_2570; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2572 = 8'hc == io_in_2 ? 8'h48 : _GEN_2571; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2573 = 8'hd == io_in_2 ? 8'h46 : _GEN_2572; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2574 = 8'he == io_in_2 ? 8'h54 : _GEN_2573; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2575 = 8'hf == io_in_2 ? 8'h5a : _GEN_2574; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2576 = 8'h10 == io_in_2 ? 8'he0 : _GEN_2575; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2577 = 8'h11 == io_in_2 ? 8'hee : _GEN_2576; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2578 = 8'h12 == io_in_2 ? 8'hfc : _GEN_2577; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2579 = 8'h13 == io_in_2 ? 8'hf2 : _GEN_2578; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2580 = 8'h14 == io_in_2 ? 8'hd8 : _GEN_2579; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2581 = 8'h15 == io_in_2 ? 8'hd6 : _GEN_2580; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2582 = 8'h16 == io_in_2 ? 8'hc4 : _GEN_2581; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2583 = 8'h17 == io_in_2 ? 8'hca : _GEN_2582; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2584 = 8'h18 == io_in_2 ? 8'h90 : _GEN_2583; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2585 = 8'h19 == io_in_2 ? 8'h9e : _GEN_2584; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2586 = 8'h1a == io_in_2 ? 8'h8c : _GEN_2585; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2587 = 8'h1b == io_in_2 ? 8'h82 : _GEN_2586; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2588 = 8'h1c == io_in_2 ? 8'ha8 : _GEN_2587; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2589 = 8'h1d == io_in_2 ? 8'ha6 : _GEN_2588; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2590 = 8'h1e == io_in_2 ? 8'hb4 : _GEN_2589; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2591 = 8'h1f == io_in_2 ? 8'hba : _GEN_2590; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2592 = 8'h20 == io_in_2 ? 8'hdb : _GEN_2591; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2593 = 8'h21 == io_in_2 ? 8'hd5 : _GEN_2592; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2594 = 8'h22 == io_in_2 ? 8'hc7 : _GEN_2593; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2595 = 8'h23 == io_in_2 ? 8'hc9 : _GEN_2594; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2596 = 8'h24 == io_in_2 ? 8'he3 : _GEN_2595; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2597 = 8'h25 == io_in_2 ? 8'hed : _GEN_2596; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2598 = 8'h26 == io_in_2 ? 8'hff : _GEN_2597; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2599 = 8'h27 == io_in_2 ? 8'hf1 : _GEN_2598; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2600 = 8'h28 == io_in_2 ? 8'hab : _GEN_2599; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2601 = 8'h29 == io_in_2 ? 8'ha5 : _GEN_2600; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2602 = 8'h2a == io_in_2 ? 8'hb7 : _GEN_2601; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2603 = 8'h2b == io_in_2 ? 8'hb9 : _GEN_2602; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2604 = 8'h2c == io_in_2 ? 8'h93 : _GEN_2603; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2605 = 8'h2d == io_in_2 ? 8'h9d : _GEN_2604; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2606 = 8'h2e == io_in_2 ? 8'h8f : _GEN_2605; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2607 = 8'h2f == io_in_2 ? 8'h81 : _GEN_2606; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2608 = 8'h30 == io_in_2 ? 8'h3b : _GEN_2607; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2609 = 8'h31 == io_in_2 ? 8'h35 : _GEN_2608; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2610 = 8'h32 == io_in_2 ? 8'h27 : _GEN_2609; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2611 = 8'h33 == io_in_2 ? 8'h29 : _GEN_2610; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2612 = 8'h34 == io_in_2 ? 8'h3 : _GEN_2611; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2613 = 8'h35 == io_in_2 ? 8'hd : _GEN_2612; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2614 = 8'h36 == io_in_2 ? 8'h1f : _GEN_2613; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2615 = 8'h37 == io_in_2 ? 8'h11 : _GEN_2614; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2616 = 8'h38 == io_in_2 ? 8'h4b : _GEN_2615; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2617 = 8'h39 == io_in_2 ? 8'h45 : _GEN_2616; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2618 = 8'h3a == io_in_2 ? 8'h57 : _GEN_2617; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2619 = 8'h3b == io_in_2 ? 8'h59 : _GEN_2618; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2620 = 8'h3c == io_in_2 ? 8'h73 : _GEN_2619; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2621 = 8'h3d == io_in_2 ? 8'h7d : _GEN_2620; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2622 = 8'h3e == io_in_2 ? 8'h6f : _GEN_2621; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2623 = 8'h3f == io_in_2 ? 8'h61 : _GEN_2622; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2624 = 8'h40 == io_in_2 ? 8'had : _GEN_2623; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2625 = 8'h41 == io_in_2 ? 8'ha3 : _GEN_2624; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2626 = 8'h42 == io_in_2 ? 8'hb1 : _GEN_2625; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2627 = 8'h43 == io_in_2 ? 8'hbf : _GEN_2626; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2628 = 8'h44 == io_in_2 ? 8'h95 : _GEN_2627; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2629 = 8'h45 == io_in_2 ? 8'h9b : _GEN_2628; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2630 = 8'h46 == io_in_2 ? 8'h89 : _GEN_2629; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2631 = 8'h47 == io_in_2 ? 8'h87 : _GEN_2630; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2632 = 8'h48 == io_in_2 ? 8'hdd : _GEN_2631; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2633 = 8'h49 == io_in_2 ? 8'hd3 : _GEN_2632; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2634 = 8'h4a == io_in_2 ? 8'hc1 : _GEN_2633; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2635 = 8'h4b == io_in_2 ? 8'hcf : _GEN_2634; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2636 = 8'h4c == io_in_2 ? 8'he5 : _GEN_2635; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2637 = 8'h4d == io_in_2 ? 8'heb : _GEN_2636; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2638 = 8'h4e == io_in_2 ? 8'hf9 : _GEN_2637; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2639 = 8'h4f == io_in_2 ? 8'hf7 : _GEN_2638; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2640 = 8'h50 == io_in_2 ? 8'h4d : _GEN_2639; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2641 = 8'h51 == io_in_2 ? 8'h43 : _GEN_2640; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2642 = 8'h52 == io_in_2 ? 8'h51 : _GEN_2641; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2643 = 8'h53 == io_in_2 ? 8'h5f : _GEN_2642; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2644 = 8'h54 == io_in_2 ? 8'h75 : _GEN_2643; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2645 = 8'h55 == io_in_2 ? 8'h7b : _GEN_2644; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2646 = 8'h56 == io_in_2 ? 8'h69 : _GEN_2645; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2647 = 8'h57 == io_in_2 ? 8'h67 : _GEN_2646; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2648 = 8'h58 == io_in_2 ? 8'h3d : _GEN_2647; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2649 = 8'h59 == io_in_2 ? 8'h33 : _GEN_2648; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2650 = 8'h5a == io_in_2 ? 8'h21 : _GEN_2649; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2651 = 8'h5b == io_in_2 ? 8'h2f : _GEN_2650; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2652 = 8'h5c == io_in_2 ? 8'h5 : _GEN_2651; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2653 = 8'h5d == io_in_2 ? 8'hb : _GEN_2652; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2654 = 8'h5e == io_in_2 ? 8'h19 : _GEN_2653; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2655 = 8'h5f == io_in_2 ? 8'h17 : _GEN_2654; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2656 = 8'h60 == io_in_2 ? 8'h76 : _GEN_2655; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2657 = 8'h61 == io_in_2 ? 8'h78 : _GEN_2656; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2658 = 8'h62 == io_in_2 ? 8'h6a : _GEN_2657; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2659 = 8'h63 == io_in_2 ? 8'h64 : _GEN_2658; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2660 = 8'h64 == io_in_2 ? 8'h4e : _GEN_2659; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2661 = 8'h65 == io_in_2 ? 8'h40 : _GEN_2660; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2662 = 8'h66 == io_in_2 ? 8'h52 : _GEN_2661; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2663 = 8'h67 == io_in_2 ? 8'h5c : _GEN_2662; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2664 = 8'h68 == io_in_2 ? 8'h6 : _GEN_2663; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2665 = 8'h69 == io_in_2 ? 8'h8 : _GEN_2664; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2666 = 8'h6a == io_in_2 ? 8'h1a : _GEN_2665; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2667 = 8'h6b == io_in_2 ? 8'h14 : _GEN_2666; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2668 = 8'h6c == io_in_2 ? 8'h3e : _GEN_2667; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2669 = 8'h6d == io_in_2 ? 8'h30 : _GEN_2668; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2670 = 8'h6e == io_in_2 ? 8'h22 : _GEN_2669; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2671 = 8'h6f == io_in_2 ? 8'h2c : _GEN_2670; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2672 = 8'h70 == io_in_2 ? 8'h96 : _GEN_2671; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2673 = 8'h71 == io_in_2 ? 8'h98 : _GEN_2672; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2674 = 8'h72 == io_in_2 ? 8'h8a : _GEN_2673; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2675 = 8'h73 == io_in_2 ? 8'h84 : _GEN_2674; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2676 = 8'h74 == io_in_2 ? 8'hae : _GEN_2675; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2677 = 8'h75 == io_in_2 ? 8'ha0 : _GEN_2676; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2678 = 8'h76 == io_in_2 ? 8'hb2 : _GEN_2677; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2679 = 8'h77 == io_in_2 ? 8'hbc : _GEN_2678; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2680 = 8'h78 == io_in_2 ? 8'he6 : _GEN_2679; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2681 = 8'h79 == io_in_2 ? 8'he8 : _GEN_2680; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2682 = 8'h7a == io_in_2 ? 8'hfa : _GEN_2681; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2683 = 8'h7b == io_in_2 ? 8'hf4 : _GEN_2682; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2684 = 8'h7c == io_in_2 ? 8'hde : _GEN_2683; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2685 = 8'h7d == io_in_2 ? 8'hd0 : _GEN_2684; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2686 = 8'h7e == io_in_2 ? 8'hc2 : _GEN_2685; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2687 = 8'h7f == io_in_2 ? 8'hcc : _GEN_2686; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2688 = 8'h80 == io_in_2 ? 8'h41 : _GEN_2687; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2689 = 8'h81 == io_in_2 ? 8'h4f : _GEN_2688; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2690 = 8'h82 == io_in_2 ? 8'h5d : _GEN_2689; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2691 = 8'h83 == io_in_2 ? 8'h53 : _GEN_2690; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2692 = 8'h84 == io_in_2 ? 8'h79 : _GEN_2691; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2693 = 8'h85 == io_in_2 ? 8'h77 : _GEN_2692; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2694 = 8'h86 == io_in_2 ? 8'h65 : _GEN_2693; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2695 = 8'h87 == io_in_2 ? 8'h6b : _GEN_2694; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2696 = 8'h88 == io_in_2 ? 8'h31 : _GEN_2695; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2697 = 8'h89 == io_in_2 ? 8'h3f : _GEN_2696; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2698 = 8'h8a == io_in_2 ? 8'h2d : _GEN_2697; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2699 = 8'h8b == io_in_2 ? 8'h23 : _GEN_2698; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2700 = 8'h8c == io_in_2 ? 8'h9 : _GEN_2699; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2701 = 8'h8d == io_in_2 ? 8'h7 : _GEN_2700; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2702 = 8'h8e == io_in_2 ? 8'h15 : _GEN_2701; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2703 = 8'h8f == io_in_2 ? 8'h1b : _GEN_2702; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2704 = 8'h90 == io_in_2 ? 8'ha1 : _GEN_2703; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2705 = 8'h91 == io_in_2 ? 8'haf : _GEN_2704; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2706 = 8'h92 == io_in_2 ? 8'hbd : _GEN_2705; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2707 = 8'h93 == io_in_2 ? 8'hb3 : _GEN_2706; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2708 = 8'h94 == io_in_2 ? 8'h99 : _GEN_2707; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2709 = 8'h95 == io_in_2 ? 8'h97 : _GEN_2708; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2710 = 8'h96 == io_in_2 ? 8'h85 : _GEN_2709; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2711 = 8'h97 == io_in_2 ? 8'h8b : _GEN_2710; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2712 = 8'h98 == io_in_2 ? 8'hd1 : _GEN_2711; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2713 = 8'h99 == io_in_2 ? 8'hdf : _GEN_2712; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2714 = 8'h9a == io_in_2 ? 8'hcd : _GEN_2713; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2715 = 8'h9b == io_in_2 ? 8'hc3 : _GEN_2714; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2716 = 8'h9c == io_in_2 ? 8'he9 : _GEN_2715; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2717 = 8'h9d == io_in_2 ? 8'he7 : _GEN_2716; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2718 = 8'h9e == io_in_2 ? 8'hf5 : _GEN_2717; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2719 = 8'h9f == io_in_2 ? 8'hfb : _GEN_2718; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2720 = 8'ha0 == io_in_2 ? 8'h9a : _GEN_2719; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2721 = 8'ha1 == io_in_2 ? 8'h94 : _GEN_2720; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2722 = 8'ha2 == io_in_2 ? 8'h86 : _GEN_2721; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2723 = 8'ha3 == io_in_2 ? 8'h88 : _GEN_2722; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2724 = 8'ha4 == io_in_2 ? 8'ha2 : _GEN_2723; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2725 = 8'ha5 == io_in_2 ? 8'hac : _GEN_2724; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2726 = 8'ha6 == io_in_2 ? 8'hbe : _GEN_2725; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2727 = 8'ha7 == io_in_2 ? 8'hb0 : _GEN_2726; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2728 = 8'ha8 == io_in_2 ? 8'hea : _GEN_2727; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2729 = 8'ha9 == io_in_2 ? 8'he4 : _GEN_2728; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2730 = 8'haa == io_in_2 ? 8'hf6 : _GEN_2729; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2731 = 8'hab == io_in_2 ? 8'hf8 : _GEN_2730; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2732 = 8'hac == io_in_2 ? 8'hd2 : _GEN_2731; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2733 = 8'had == io_in_2 ? 8'hdc : _GEN_2732; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2734 = 8'hae == io_in_2 ? 8'hce : _GEN_2733; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2735 = 8'haf == io_in_2 ? 8'hc0 : _GEN_2734; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2736 = 8'hb0 == io_in_2 ? 8'h7a : _GEN_2735; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2737 = 8'hb1 == io_in_2 ? 8'h74 : _GEN_2736; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2738 = 8'hb2 == io_in_2 ? 8'h66 : _GEN_2737; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2739 = 8'hb3 == io_in_2 ? 8'h68 : _GEN_2738; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2740 = 8'hb4 == io_in_2 ? 8'h42 : _GEN_2739; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2741 = 8'hb5 == io_in_2 ? 8'h4c : _GEN_2740; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2742 = 8'hb6 == io_in_2 ? 8'h5e : _GEN_2741; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2743 = 8'hb7 == io_in_2 ? 8'h50 : _GEN_2742; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2744 = 8'hb8 == io_in_2 ? 8'ha : _GEN_2743; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2745 = 8'hb9 == io_in_2 ? 8'h4 : _GEN_2744; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2746 = 8'hba == io_in_2 ? 8'h16 : _GEN_2745; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2747 = 8'hbb == io_in_2 ? 8'h18 : _GEN_2746; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2748 = 8'hbc == io_in_2 ? 8'h32 : _GEN_2747; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2749 = 8'hbd == io_in_2 ? 8'h3c : _GEN_2748; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2750 = 8'hbe == io_in_2 ? 8'h2e : _GEN_2749; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2751 = 8'hbf == io_in_2 ? 8'h20 : _GEN_2750; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2752 = 8'hc0 == io_in_2 ? 8'hec : _GEN_2751; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2753 = 8'hc1 == io_in_2 ? 8'he2 : _GEN_2752; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2754 = 8'hc2 == io_in_2 ? 8'hf0 : _GEN_2753; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2755 = 8'hc3 == io_in_2 ? 8'hfe : _GEN_2754; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2756 = 8'hc4 == io_in_2 ? 8'hd4 : _GEN_2755; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2757 = 8'hc5 == io_in_2 ? 8'hda : _GEN_2756; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2758 = 8'hc6 == io_in_2 ? 8'hc8 : _GEN_2757; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2759 = 8'hc7 == io_in_2 ? 8'hc6 : _GEN_2758; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2760 = 8'hc8 == io_in_2 ? 8'h9c : _GEN_2759; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2761 = 8'hc9 == io_in_2 ? 8'h92 : _GEN_2760; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2762 = 8'hca == io_in_2 ? 8'h80 : _GEN_2761; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2763 = 8'hcb == io_in_2 ? 8'h8e : _GEN_2762; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2764 = 8'hcc == io_in_2 ? 8'ha4 : _GEN_2763; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2765 = 8'hcd == io_in_2 ? 8'haa : _GEN_2764; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2766 = 8'hce == io_in_2 ? 8'hb8 : _GEN_2765; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2767 = 8'hcf == io_in_2 ? 8'hb6 : _GEN_2766; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2768 = 8'hd0 == io_in_2 ? 8'hc : _GEN_2767; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2769 = 8'hd1 == io_in_2 ? 8'h2 : _GEN_2768; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2770 = 8'hd2 == io_in_2 ? 8'h10 : _GEN_2769; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2771 = 8'hd3 == io_in_2 ? 8'h1e : _GEN_2770; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2772 = 8'hd4 == io_in_2 ? 8'h34 : _GEN_2771; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2773 = 8'hd5 == io_in_2 ? 8'h3a : _GEN_2772; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2774 = 8'hd6 == io_in_2 ? 8'h28 : _GEN_2773; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2775 = 8'hd7 == io_in_2 ? 8'h26 : _GEN_2774; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2776 = 8'hd8 == io_in_2 ? 8'h7c : _GEN_2775; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2777 = 8'hd9 == io_in_2 ? 8'h72 : _GEN_2776; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2778 = 8'hda == io_in_2 ? 8'h60 : _GEN_2777; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2779 = 8'hdb == io_in_2 ? 8'h6e : _GEN_2778; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2780 = 8'hdc == io_in_2 ? 8'h44 : _GEN_2779; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2781 = 8'hdd == io_in_2 ? 8'h4a : _GEN_2780; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2782 = 8'hde == io_in_2 ? 8'h58 : _GEN_2781; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2783 = 8'hdf == io_in_2 ? 8'h56 : _GEN_2782; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2784 = 8'he0 == io_in_2 ? 8'h37 : _GEN_2783; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2785 = 8'he1 == io_in_2 ? 8'h39 : _GEN_2784; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2786 = 8'he2 == io_in_2 ? 8'h2b : _GEN_2785; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2787 = 8'he3 == io_in_2 ? 8'h25 : _GEN_2786; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2788 = 8'he4 == io_in_2 ? 8'hf : _GEN_2787; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2789 = 8'he5 == io_in_2 ? 8'h1 : _GEN_2788; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2790 = 8'he6 == io_in_2 ? 8'h13 : _GEN_2789; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2791 = 8'he7 == io_in_2 ? 8'h1d : _GEN_2790; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2792 = 8'he8 == io_in_2 ? 8'h47 : _GEN_2791; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2793 = 8'he9 == io_in_2 ? 8'h49 : _GEN_2792; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2794 = 8'hea == io_in_2 ? 8'h5b : _GEN_2793; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2795 = 8'heb == io_in_2 ? 8'h55 : _GEN_2794; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2796 = 8'hec == io_in_2 ? 8'h7f : _GEN_2795; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2797 = 8'hed == io_in_2 ? 8'h71 : _GEN_2796; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2798 = 8'hee == io_in_2 ? 8'h63 : _GEN_2797; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2799 = 8'hef == io_in_2 ? 8'h6d : _GEN_2798; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2800 = 8'hf0 == io_in_2 ? 8'hd7 : _GEN_2799; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2801 = 8'hf1 == io_in_2 ? 8'hd9 : _GEN_2800; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2802 = 8'hf2 == io_in_2 ? 8'hcb : _GEN_2801; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2803 = 8'hf3 == io_in_2 ? 8'hc5 : _GEN_2802; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2804 = 8'hf4 == io_in_2 ? 8'hef : _GEN_2803; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2805 = 8'hf5 == io_in_2 ? 8'he1 : _GEN_2804; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2806 = 8'hf6 == io_in_2 ? 8'hf3 : _GEN_2805; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2807 = 8'hf7 == io_in_2 ? 8'hfd : _GEN_2806; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2808 = 8'hf8 == io_in_2 ? 8'ha7 : _GEN_2807; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2809 = 8'hf9 == io_in_2 ? 8'ha9 : _GEN_2808; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2810 = 8'hfa == io_in_2 ? 8'hbb : _GEN_2809; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2811 = 8'hfb == io_in_2 ? 8'hb5 : _GEN_2810; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2812 = 8'hfc == io_in_2 ? 8'h9f : _GEN_2811; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2813 = 8'hfd == io_in_2 ? 8'h91 : _GEN_2812; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2814 = 8'hfe == io_in_2 ? 8'h83 : _GEN_2813; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2815 = 8'hff == io_in_2 ? 8'h8d : _GEN_2814; // @[AES_PipelinedElasticBuffer.scala 593:49 AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _T_7 = _T_6 ^ _GEN_2815; // @[AES_PipelinedElasticBuffer.scala 593:49]
  wire [7:0] _GEN_2817 = 8'h1 == io_in_3 ? 8'hb : 8'h0; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2818 = 8'h2 == io_in_3 ? 8'h16 : _GEN_2817; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2819 = 8'h3 == io_in_3 ? 8'h1d : _GEN_2818; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2820 = 8'h4 == io_in_3 ? 8'h2c : _GEN_2819; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2821 = 8'h5 == io_in_3 ? 8'h27 : _GEN_2820; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2822 = 8'h6 == io_in_3 ? 8'h3a : _GEN_2821; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2823 = 8'h7 == io_in_3 ? 8'h31 : _GEN_2822; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2824 = 8'h8 == io_in_3 ? 8'h58 : _GEN_2823; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2825 = 8'h9 == io_in_3 ? 8'h53 : _GEN_2824; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2826 = 8'ha == io_in_3 ? 8'h4e : _GEN_2825; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2827 = 8'hb == io_in_3 ? 8'h45 : _GEN_2826; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2828 = 8'hc == io_in_3 ? 8'h74 : _GEN_2827; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2829 = 8'hd == io_in_3 ? 8'h7f : _GEN_2828; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2830 = 8'he == io_in_3 ? 8'h62 : _GEN_2829; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2831 = 8'hf == io_in_3 ? 8'h69 : _GEN_2830; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2832 = 8'h10 == io_in_3 ? 8'hb0 : _GEN_2831; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2833 = 8'h11 == io_in_3 ? 8'hbb : _GEN_2832; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2834 = 8'h12 == io_in_3 ? 8'ha6 : _GEN_2833; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2835 = 8'h13 == io_in_3 ? 8'had : _GEN_2834; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2836 = 8'h14 == io_in_3 ? 8'h9c : _GEN_2835; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2837 = 8'h15 == io_in_3 ? 8'h97 : _GEN_2836; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2838 = 8'h16 == io_in_3 ? 8'h8a : _GEN_2837; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2839 = 8'h17 == io_in_3 ? 8'h81 : _GEN_2838; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2840 = 8'h18 == io_in_3 ? 8'he8 : _GEN_2839; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2841 = 8'h19 == io_in_3 ? 8'he3 : _GEN_2840; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2842 = 8'h1a == io_in_3 ? 8'hfe : _GEN_2841; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2843 = 8'h1b == io_in_3 ? 8'hf5 : _GEN_2842; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2844 = 8'h1c == io_in_3 ? 8'hc4 : _GEN_2843; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2845 = 8'h1d == io_in_3 ? 8'hcf : _GEN_2844; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2846 = 8'h1e == io_in_3 ? 8'hd2 : _GEN_2845; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2847 = 8'h1f == io_in_3 ? 8'hd9 : _GEN_2846; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2848 = 8'h20 == io_in_3 ? 8'h7b : _GEN_2847; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2849 = 8'h21 == io_in_3 ? 8'h70 : _GEN_2848; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2850 = 8'h22 == io_in_3 ? 8'h6d : _GEN_2849; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2851 = 8'h23 == io_in_3 ? 8'h66 : _GEN_2850; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2852 = 8'h24 == io_in_3 ? 8'h57 : _GEN_2851; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2853 = 8'h25 == io_in_3 ? 8'h5c : _GEN_2852; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2854 = 8'h26 == io_in_3 ? 8'h41 : _GEN_2853; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2855 = 8'h27 == io_in_3 ? 8'h4a : _GEN_2854; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2856 = 8'h28 == io_in_3 ? 8'h23 : _GEN_2855; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2857 = 8'h29 == io_in_3 ? 8'h28 : _GEN_2856; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2858 = 8'h2a == io_in_3 ? 8'h35 : _GEN_2857; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2859 = 8'h2b == io_in_3 ? 8'h3e : _GEN_2858; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2860 = 8'h2c == io_in_3 ? 8'hf : _GEN_2859; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2861 = 8'h2d == io_in_3 ? 8'h4 : _GEN_2860; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2862 = 8'h2e == io_in_3 ? 8'h19 : _GEN_2861; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2863 = 8'h2f == io_in_3 ? 8'h12 : _GEN_2862; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2864 = 8'h30 == io_in_3 ? 8'hcb : _GEN_2863; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2865 = 8'h31 == io_in_3 ? 8'hc0 : _GEN_2864; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2866 = 8'h32 == io_in_3 ? 8'hdd : _GEN_2865; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2867 = 8'h33 == io_in_3 ? 8'hd6 : _GEN_2866; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2868 = 8'h34 == io_in_3 ? 8'he7 : _GEN_2867; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2869 = 8'h35 == io_in_3 ? 8'hec : _GEN_2868; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2870 = 8'h36 == io_in_3 ? 8'hf1 : _GEN_2869; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2871 = 8'h37 == io_in_3 ? 8'hfa : _GEN_2870; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2872 = 8'h38 == io_in_3 ? 8'h93 : _GEN_2871; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2873 = 8'h39 == io_in_3 ? 8'h98 : _GEN_2872; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2874 = 8'h3a == io_in_3 ? 8'h85 : _GEN_2873; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2875 = 8'h3b == io_in_3 ? 8'h8e : _GEN_2874; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2876 = 8'h3c == io_in_3 ? 8'hbf : _GEN_2875; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2877 = 8'h3d == io_in_3 ? 8'hb4 : _GEN_2876; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2878 = 8'h3e == io_in_3 ? 8'ha9 : _GEN_2877; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2879 = 8'h3f == io_in_3 ? 8'ha2 : _GEN_2878; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2880 = 8'h40 == io_in_3 ? 8'hf6 : _GEN_2879; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2881 = 8'h41 == io_in_3 ? 8'hfd : _GEN_2880; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2882 = 8'h42 == io_in_3 ? 8'he0 : _GEN_2881; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2883 = 8'h43 == io_in_3 ? 8'heb : _GEN_2882; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2884 = 8'h44 == io_in_3 ? 8'hda : _GEN_2883; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2885 = 8'h45 == io_in_3 ? 8'hd1 : _GEN_2884; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2886 = 8'h46 == io_in_3 ? 8'hcc : _GEN_2885; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2887 = 8'h47 == io_in_3 ? 8'hc7 : _GEN_2886; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2888 = 8'h48 == io_in_3 ? 8'hae : _GEN_2887; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2889 = 8'h49 == io_in_3 ? 8'ha5 : _GEN_2888; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2890 = 8'h4a == io_in_3 ? 8'hb8 : _GEN_2889; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2891 = 8'h4b == io_in_3 ? 8'hb3 : _GEN_2890; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2892 = 8'h4c == io_in_3 ? 8'h82 : _GEN_2891; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2893 = 8'h4d == io_in_3 ? 8'h89 : _GEN_2892; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2894 = 8'h4e == io_in_3 ? 8'h94 : _GEN_2893; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2895 = 8'h4f == io_in_3 ? 8'h9f : _GEN_2894; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2896 = 8'h50 == io_in_3 ? 8'h46 : _GEN_2895; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2897 = 8'h51 == io_in_3 ? 8'h4d : _GEN_2896; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2898 = 8'h52 == io_in_3 ? 8'h50 : _GEN_2897; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2899 = 8'h53 == io_in_3 ? 8'h5b : _GEN_2898; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2900 = 8'h54 == io_in_3 ? 8'h6a : _GEN_2899; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2901 = 8'h55 == io_in_3 ? 8'h61 : _GEN_2900; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2902 = 8'h56 == io_in_3 ? 8'h7c : _GEN_2901; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2903 = 8'h57 == io_in_3 ? 8'h77 : _GEN_2902; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2904 = 8'h58 == io_in_3 ? 8'h1e : _GEN_2903; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2905 = 8'h59 == io_in_3 ? 8'h15 : _GEN_2904; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2906 = 8'h5a == io_in_3 ? 8'h8 : _GEN_2905; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2907 = 8'h5b == io_in_3 ? 8'h3 : _GEN_2906; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2908 = 8'h5c == io_in_3 ? 8'h32 : _GEN_2907; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2909 = 8'h5d == io_in_3 ? 8'h39 : _GEN_2908; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2910 = 8'h5e == io_in_3 ? 8'h24 : _GEN_2909; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2911 = 8'h5f == io_in_3 ? 8'h2f : _GEN_2910; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2912 = 8'h60 == io_in_3 ? 8'h8d : _GEN_2911; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2913 = 8'h61 == io_in_3 ? 8'h86 : _GEN_2912; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2914 = 8'h62 == io_in_3 ? 8'h9b : _GEN_2913; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2915 = 8'h63 == io_in_3 ? 8'h90 : _GEN_2914; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2916 = 8'h64 == io_in_3 ? 8'ha1 : _GEN_2915; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2917 = 8'h65 == io_in_3 ? 8'haa : _GEN_2916; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2918 = 8'h66 == io_in_3 ? 8'hb7 : _GEN_2917; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2919 = 8'h67 == io_in_3 ? 8'hbc : _GEN_2918; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2920 = 8'h68 == io_in_3 ? 8'hd5 : _GEN_2919; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2921 = 8'h69 == io_in_3 ? 8'hde : _GEN_2920; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2922 = 8'h6a == io_in_3 ? 8'hc3 : _GEN_2921; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2923 = 8'h6b == io_in_3 ? 8'hc8 : _GEN_2922; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2924 = 8'h6c == io_in_3 ? 8'hf9 : _GEN_2923; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2925 = 8'h6d == io_in_3 ? 8'hf2 : _GEN_2924; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2926 = 8'h6e == io_in_3 ? 8'hef : _GEN_2925; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2927 = 8'h6f == io_in_3 ? 8'he4 : _GEN_2926; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2928 = 8'h70 == io_in_3 ? 8'h3d : _GEN_2927; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2929 = 8'h71 == io_in_3 ? 8'h36 : _GEN_2928; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2930 = 8'h72 == io_in_3 ? 8'h2b : _GEN_2929; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2931 = 8'h73 == io_in_3 ? 8'h20 : _GEN_2930; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2932 = 8'h74 == io_in_3 ? 8'h11 : _GEN_2931; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2933 = 8'h75 == io_in_3 ? 8'h1a : _GEN_2932; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2934 = 8'h76 == io_in_3 ? 8'h7 : _GEN_2933; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2935 = 8'h77 == io_in_3 ? 8'hc : _GEN_2934; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2936 = 8'h78 == io_in_3 ? 8'h65 : _GEN_2935; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2937 = 8'h79 == io_in_3 ? 8'h6e : _GEN_2936; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2938 = 8'h7a == io_in_3 ? 8'h73 : _GEN_2937; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2939 = 8'h7b == io_in_3 ? 8'h78 : _GEN_2938; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2940 = 8'h7c == io_in_3 ? 8'h49 : _GEN_2939; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2941 = 8'h7d == io_in_3 ? 8'h42 : _GEN_2940; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2942 = 8'h7e == io_in_3 ? 8'h5f : _GEN_2941; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2943 = 8'h7f == io_in_3 ? 8'h54 : _GEN_2942; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2944 = 8'h80 == io_in_3 ? 8'hf7 : _GEN_2943; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2945 = 8'h81 == io_in_3 ? 8'hfc : _GEN_2944; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2946 = 8'h82 == io_in_3 ? 8'he1 : _GEN_2945; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2947 = 8'h83 == io_in_3 ? 8'hea : _GEN_2946; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2948 = 8'h84 == io_in_3 ? 8'hdb : _GEN_2947; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2949 = 8'h85 == io_in_3 ? 8'hd0 : _GEN_2948; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2950 = 8'h86 == io_in_3 ? 8'hcd : _GEN_2949; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2951 = 8'h87 == io_in_3 ? 8'hc6 : _GEN_2950; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2952 = 8'h88 == io_in_3 ? 8'haf : _GEN_2951; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2953 = 8'h89 == io_in_3 ? 8'ha4 : _GEN_2952; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2954 = 8'h8a == io_in_3 ? 8'hb9 : _GEN_2953; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2955 = 8'h8b == io_in_3 ? 8'hb2 : _GEN_2954; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2956 = 8'h8c == io_in_3 ? 8'h83 : _GEN_2955; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2957 = 8'h8d == io_in_3 ? 8'h88 : _GEN_2956; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2958 = 8'h8e == io_in_3 ? 8'h95 : _GEN_2957; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2959 = 8'h8f == io_in_3 ? 8'h9e : _GEN_2958; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2960 = 8'h90 == io_in_3 ? 8'h47 : _GEN_2959; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2961 = 8'h91 == io_in_3 ? 8'h4c : _GEN_2960; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2962 = 8'h92 == io_in_3 ? 8'h51 : _GEN_2961; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2963 = 8'h93 == io_in_3 ? 8'h5a : _GEN_2962; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2964 = 8'h94 == io_in_3 ? 8'h6b : _GEN_2963; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2965 = 8'h95 == io_in_3 ? 8'h60 : _GEN_2964; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2966 = 8'h96 == io_in_3 ? 8'h7d : _GEN_2965; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2967 = 8'h97 == io_in_3 ? 8'h76 : _GEN_2966; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2968 = 8'h98 == io_in_3 ? 8'h1f : _GEN_2967; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2969 = 8'h99 == io_in_3 ? 8'h14 : _GEN_2968; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2970 = 8'h9a == io_in_3 ? 8'h9 : _GEN_2969; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2971 = 8'h9b == io_in_3 ? 8'h2 : _GEN_2970; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2972 = 8'h9c == io_in_3 ? 8'h33 : _GEN_2971; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2973 = 8'h9d == io_in_3 ? 8'h38 : _GEN_2972; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2974 = 8'h9e == io_in_3 ? 8'h25 : _GEN_2973; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2975 = 8'h9f == io_in_3 ? 8'h2e : _GEN_2974; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2976 = 8'ha0 == io_in_3 ? 8'h8c : _GEN_2975; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2977 = 8'ha1 == io_in_3 ? 8'h87 : _GEN_2976; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2978 = 8'ha2 == io_in_3 ? 8'h9a : _GEN_2977; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2979 = 8'ha3 == io_in_3 ? 8'h91 : _GEN_2978; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2980 = 8'ha4 == io_in_3 ? 8'ha0 : _GEN_2979; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2981 = 8'ha5 == io_in_3 ? 8'hab : _GEN_2980; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2982 = 8'ha6 == io_in_3 ? 8'hb6 : _GEN_2981; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2983 = 8'ha7 == io_in_3 ? 8'hbd : _GEN_2982; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2984 = 8'ha8 == io_in_3 ? 8'hd4 : _GEN_2983; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2985 = 8'ha9 == io_in_3 ? 8'hdf : _GEN_2984; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2986 = 8'haa == io_in_3 ? 8'hc2 : _GEN_2985; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2987 = 8'hab == io_in_3 ? 8'hc9 : _GEN_2986; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2988 = 8'hac == io_in_3 ? 8'hf8 : _GEN_2987; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2989 = 8'had == io_in_3 ? 8'hf3 : _GEN_2988; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2990 = 8'hae == io_in_3 ? 8'hee : _GEN_2989; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2991 = 8'haf == io_in_3 ? 8'he5 : _GEN_2990; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2992 = 8'hb0 == io_in_3 ? 8'h3c : _GEN_2991; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2993 = 8'hb1 == io_in_3 ? 8'h37 : _GEN_2992; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2994 = 8'hb2 == io_in_3 ? 8'h2a : _GEN_2993; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2995 = 8'hb3 == io_in_3 ? 8'h21 : _GEN_2994; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2996 = 8'hb4 == io_in_3 ? 8'h10 : _GEN_2995; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2997 = 8'hb5 == io_in_3 ? 8'h1b : _GEN_2996; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2998 = 8'hb6 == io_in_3 ? 8'h6 : _GEN_2997; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_2999 = 8'hb7 == io_in_3 ? 8'hd : _GEN_2998; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3000 = 8'hb8 == io_in_3 ? 8'h64 : _GEN_2999; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3001 = 8'hb9 == io_in_3 ? 8'h6f : _GEN_3000; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3002 = 8'hba == io_in_3 ? 8'h72 : _GEN_3001; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3003 = 8'hbb == io_in_3 ? 8'h79 : _GEN_3002; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3004 = 8'hbc == io_in_3 ? 8'h48 : _GEN_3003; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3005 = 8'hbd == io_in_3 ? 8'h43 : _GEN_3004; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3006 = 8'hbe == io_in_3 ? 8'h5e : _GEN_3005; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3007 = 8'hbf == io_in_3 ? 8'h55 : _GEN_3006; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3008 = 8'hc0 == io_in_3 ? 8'h1 : _GEN_3007; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3009 = 8'hc1 == io_in_3 ? 8'ha : _GEN_3008; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3010 = 8'hc2 == io_in_3 ? 8'h17 : _GEN_3009; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3011 = 8'hc3 == io_in_3 ? 8'h1c : _GEN_3010; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3012 = 8'hc4 == io_in_3 ? 8'h2d : _GEN_3011; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3013 = 8'hc5 == io_in_3 ? 8'h26 : _GEN_3012; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3014 = 8'hc6 == io_in_3 ? 8'h3b : _GEN_3013; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3015 = 8'hc7 == io_in_3 ? 8'h30 : _GEN_3014; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3016 = 8'hc8 == io_in_3 ? 8'h59 : _GEN_3015; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3017 = 8'hc9 == io_in_3 ? 8'h52 : _GEN_3016; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3018 = 8'hca == io_in_3 ? 8'h4f : _GEN_3017; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3019 = 8'hcb == io_in_3 ? 8'h44 : _GEN_3018; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3020 = 8'hcc == io_in_3 ? 8'h75 : _GEN_3019; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3021 = 8'hcd == io_in_3 ? 8'h7e : _GEN_3020; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3022 = 8'hce == io_in_3 ? 8'h63 : _GEN_3021; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3023 = 8'hcf == io_in_3 ? 8'h68 : _GEN_3022; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3024 = 8'hd0 == io_in_3 ? 8'hb1 : _GEN_3023; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3025 = 8'hd1 == io_in_3 ? 8'hba : _GEN_3024; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3026 = 8'hd2 == io_in_3 ? 8'ha7 : _GEN_3025; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3027 = 8'hd3 == io_in_3 ? 8'hac : _GEN_3026; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3028 = 8'hd4 == io_in_3 ? 8'h9d : _GEN_3027; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3029 = 8'hd5 == io_in_3 ? 8'h96 : _GEN_3028; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3030 = 8'hd6 == io_in_3 ? 8'h8b : _GEN_3029; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3031 = 8'hd7 == io_in_3 ? 8'h80 : _GEN_3030; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3032 = 8'hd8 == io_in_3 ? 8'he9 : _GEN_3031; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3033 = 8'hd9 == io_in_3 ? 8'he2 : _GEN_3032; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3034 = 8'hda == io_in_3 ? 8'hff : _GEN_3033; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3035 = 8'hdb == io_in_3 ? 8'hf4 : _GEN_3034; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3036 = 8'hdc == io_in_3 ? 8'hc5 : _GEN_3035; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3037 = 8'hdd == io_in_3 ? 8'hce : _GEN_3036; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3038 = 8'hde == io_in_3 ? 8'hd3 : _GEN_3037; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3039 = 8'hdf == io_in_3 ? 8'hd8 : _GEN_3038; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3040 = 8'he0 == io_in_3 ? 8'h7a : _GEN_3039; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3041 = 8'he1 == io_in_3 ? 8'h71 : _GEN_3040; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3042 = 8'he2 == io_in_3 ? 8'h6c : _GEN_3041; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3043 = 8'he3 == io_in_3 ? 8'h67 : _GEN_3042; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3044 = 8'he4 == io_in_3 ? 8'h56 : _GEN_3043; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3045 = 8'he5 == io_in_3 ? 8'h5d : _GEN_3044; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3046 = 8'he6 == io_in_3 ? 8'h40 : _GEN_3045; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3047 = 8'he7 == io_in_3 ? 8'h4b : _GEN_3046; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3048 = 8'he8 == io_in_3 ? 8'h22 : _GEN_3047; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3049 = 8'he9 == io_in_3 ? 8'h29 : _GEN_3048; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3050 = 8'hea == io_in_3 ? 8'h34 : _GEN_3049; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3051 = 8'heb == io_in_3 ? 8'h3f : _GEN_3050; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3052 = 8'hec == io_in_3 ? 8'he : _GEN_3051; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3053 = 8'hed == io_in_3 ? 8'h5 : _GEN_3052; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3054 = 8'hee == io_in_3 ? 8'h18 : _GEN_3053; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3055 = 8'hef == io_in_3 ? 8'h13 : _GEN_3054; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3056 = 8'hf0 == io_in_3 ? 8'hca : _GEN_3055; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3057 = 8'hf1 == io_in_3 ? 8'hc1 : _GEN_3056; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3058 = 8'hf2 == io_in_3 ? 8'hdc : _GEN_3057; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3059 = 8'hf3 == io_in_3 ? 8'hd7 : _GEN_3058; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3060 = 8'hf4 == io_in_3 ? 8'he6 : _GEN_3059; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3061 = 8'hf5 == io_in_3 ? 8'hed : _GEN_3060; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3062 = 8'hf6 == io_in_3 ? 8'hf0 : _GEN_3061; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3063 = 8'hf7 == io_in_3 ? 8'hfb : _GEN_3062; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3064 = 8'hf8 == io_in_3 ? 8'h92 : _GEN_3063; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3065 = 8'hf9 == io_in_3 ? 8'h99 : _GEN_3064; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3066 = 8'hfa == io_in_3 ? 8'h84 : _GEN_3065; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3067 = 8'hfb == io_in_3 ? 8'h8f : _GEN_3066; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3068 = 8'hfc == io_in_3 ? 8'hbe : _GEN_3067; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3069 = 8'hfd == io_in_3 ? 8'hb5 : _GEN_3068; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3070 = 8'hfe == io_in_3 ? 8'ha8 : _GEN_3069; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3071 = 8'hff == io_in_3 ? 8'ha3 : _GEN_3070; // @[AES_PipelinedElasticBuffer.scala 593:67 AES_PipelinedElasticBuffer.scala 593:67]
  wire [7:0] _GEN_3073 = 8'h1 == io_in_0 ? 8'hb : 8'h0; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3074 = 8'h2 == io_in_0 ? 8'h16 : _GEN_3073; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3075 = 8'h3 == io_in_0 ? 8'h1d : _GEN_3074; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3076 = 8'h4 == io_in_0 ? 8'h2c : _GEN_3075; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3077 = 8'h5 == io_in_0 ? 8'h27 : _GEN_3076; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3078 = 8'h6 == io_in_0 ? 8'h3a : _GEN_3077; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3079 = 8'h7 == io_in_0 ? 8'h31 : _GEN_3078; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3080 = 8'h8 == io_in_0 ? 8'h58 : _GEN_3079; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3081 = 8'h9 == io_in_0 ? 8'h53 : _GEN_3080; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3082 = 8'ha == io_in_0 ? 8'h4e : _GEN_3081; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3083 = 8'hb == io_in_0 ? 8'h45 : _GEN_3082; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3084 = 8'hc == io_in_0 ? 8'h74 : _GEN_3083; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3085 = 8'hd == io_in_0 ? 8'h7f : _GEN_3084; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3086 = 8'he == io_in_0 ? 8'h62 : _GEN_3085; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3087 = 8'hf == io_in_0 ? 8'h69 : _GEN_3086; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3088 = 8'h10 == io_in_0 ? 8'hb0 : _GEN_3087; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3089 = 8'h11 == io_in_0 ? 8'hbb : _GEN_3088; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3090 = 8'h12 == io_in_0 ? 8'ha6 : _GEN_3089; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3091 = 8'h13 == io_in_0 ? 8'had : _GEN_3090; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3092 = 8'h14 == io_in_0 ? 8'h9c : _GEN_3091; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3093 = 8'h15 == io_in_0 ? 8'h97 : _GEN_3092; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3094 = 8'h16 == io_in_0 ? 8'h8a : _GEN_3093; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3095 = 8'h17 == io_in_0 ? 8'h81 : _GEN_3094; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3096 = 8'h18 == io_in_0 ? 8'he8 : _GEN_3095; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3097 = 8'h19 == io_in_0 ? 8'he3 : _GEN_3096; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3098 = 8'h1a == io_in_0 ? 8'hfe : _GEN_3097; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3099 = 8'h1b == io_in_0 ? 8'hf5 : _GEN_3098; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3100 = 8'h1c == io_in_0 ? 8'hc4 : _GEN_3099; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3101 = 8'h1d == io_in_0 ? 8'hcf : _GEN_3100; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3102 = 8'h1e == io_in_0 ? 8'hd2 : _GEN_3101; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3103 = 8'h1f == io_in_0 ? 8'hd9 : _GEN_3102; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3104 = 8'h20 == io_in_0 ? 8'h7b : _GEN_3103; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3105 = 8'h21 == io_in_0 ? 8'h70 : _GEN_3104; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3106 = 8'h22 == io_in_0 ? 8'h6d : _GEN_3105; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3107 = 8'h23 == io_in_0 ? 8'h66 : _GEN_3106; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3108 = 8'h24 == io_in_0 ? 8'h57 : _GEN_3107; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3109 = 8'h25 == io_in_0 ? 8'h5c : _GEN_3108; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3110 = 8'h26 == io_in_0 ? 8'h41 : _GEN_3109; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3111 = 8'h27 == io_in_0 ? 8'h4a : _GEN_3110; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3112 = 8'h28 == io_in_0 ? 8'h23 : _GEN_3111; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3113 = 8'h29 == io_in_0 ? 8'h28 : _GEN_3112; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3114 = 8'h2a == io_in_0 ? 8'h35 : _GEN_3113; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3115 = 8'h2b == io_in_0 ? 8'h3e : _GEN_3114; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3116 = 8'h2c == io_in_0 ? 8'hf : _GEN_3115; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3117 = 8'h2d == io_in_0 ? 8'h4 : _GEN_3116; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3118 = 8'h2e == io_in_0 ? 8'h19 : _GEN_3117; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3119 = 8'h2f == io_in_0 ? 8'h12 : _GEN_3118; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3120 = 8'h30 == io_in_0 ? 8'hcb : _GEN_3119; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3121 = 8'h31 == io_in_0 ? 8'hc0 : _GEN_3120; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3122 = 8'h32 == io_in_0 ? 8'hdd : _GEN_3121; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3123 = 8'h33 == io_in_0 ? 8'hd6 : _GEN_3122; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3124 = 8'h34 == io_in_0 ? 8'he7 : _GEN_3123; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3125 = 8'h35 == io_in_0 ? 8'hec : _GEN_3124; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3126 = 8'h36 == io_in_0 ? 8'hf1 : _GEN_3125; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3127 = 8'h37 == io_in_0 ? 8'hfa : _GEN_3126; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3128 = 8'h38 == io_in_0 ? 8'h93 : _GEN_3127; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3129 = 8'h39 == io_in_0 ? 8'h98 : _GEN_3128; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3130 = 8'h3a == io_in_0 ? 8'h85 : _GEN_3129; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3131 = 8'h3b == io_in_0 ? 8'h8e : _GEN_3130; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3132 = 8'h3c == io_in_0 ? 8'hbf : _GEN_3131; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3133 = 8'h3d == io_in_0 ? 8'hb4 : _GEN_3132; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3134 = 8'h3e == io_in_0 ? 8'ha9 : _GEN_3133; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3135 = 8'h3f == io_in_0 ? 8'ha2 : _GEN_3134; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3136 = 8'h40 == io_in_0 ? 8'hf6 : _GEN_3135; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3137 = 8'h41 == io_in_0 ? 8'hfd : _GEN_3136; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3138 = 8'h42 == io_in_0 ? 8'he0 : _GEN_3137; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3139 = 8'h43 == io_in_0 ? 8'heb : _GEN_3138; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3140 = 8'h44 == io_in_0 ? 8'hda : _GEN_3139; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3141 = 8'h45 == io_in_0 ? 8'hd1 : _GEN_3140; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3142 = 8'h46 == io_in_0 ? 8'hcc : _GEN_3141; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3143 = 8'h47 == io_in_0 ? 8'hc7 : _GEN_3142; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3144 = 8'h48 == io_in_0 ? 8'hae : _GEN_3143; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3145 = 8'h49 == io_in_0 ? 8'ha5 : _GEN_3144; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3146 = 8'h4a == io_in_0 ? 8'hb8 : _GEN_3145; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3147 = 8'h4b == io_in_0 ? 8'hb3 : _GEN_3146; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3148 = 8'h4c == io_in_0 ? 8'h82 : _GEN_3147; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3149 = 8'h4d == io_in_0 ? 8'h89 : _GEN_3148; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3150 = 8'h4e == io_in_0 ? 8'h94 : _GEN_3149; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3151 = 8'h4f == io_in_0 ? 8'h9f : _GEN_3150; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3152 = 8'h50 == io_in_0 ? 8'h46 : _GEN_3151; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3153 = 8'h51 == io_in_0 ? 8'h4d : _GEN_3152; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3154 = 8'h52 == io_in_0 ? 8'h50 : _GEN_3153; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3155 = 8'h53 == io_in_0 ? 8'h5b : _GEN_3154; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3156 = 8'h54 == io_in_0 ? 8'h6a : _GEN_3155; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3157 = 8'h55 == io_in_0 ? 8'h61 : _GEN_3156; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3158 = 8'h56 == io_in_0 ? 8'h7c : _GEN_3157; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3159 = 8'h57 == io_in_0 ? 8'h77 : _GEN_3158; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3160 = 8'h58 == io_in_0 ? 8'h1e : _GEN_3159; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3161 = 8'h59 == io_in_0 ? 8'h15 : _GEN_3160; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3162 = 8'h5a == io_in_0 ? 8'h8 : _GEN_3161; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3163 = 8'h5b == io_in_0 ? 8'h3 : _GEN_3162; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3164 = 8'h5c == io_in_0 ? 8'h32 : _GEN_3163; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3165 = 8'h5d == io_in_0 ? 8'h39 : _GEN_3164; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3166 = 8'h5e == io_in_0 ? 8'h24 : _GEN_3165; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3167 = 8'h5f == io_in_0 ? 8'h2f : _GEN_3166; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3168 = 8'h60 == io_in_0 ? 8'h8d : _GEN_3167; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3169 = 8'h61 == io_in_0 ? 8'h86 : _GEN_3168; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3170 = 8'h62 == io_in_0 ? 8'h9b : _GEN_3169; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3171 = 8'h63 == io_in_0 ? 8'h90 : _GEN_3170; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3172 = 8'h64 == io_in_0 ? 8'ha1 : _GEN_3171; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3173 = 8'h65 == io_in_0 ? 8'haa : _GEN_3172; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3174 = 8'h66 == io_in_0 ? 8'hb7 : _GEN_3173; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3175 = 8'h67 == io_in_0 ? 8'hbc : _GEN_3174; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3176 = 8'h68 == io_in_0 ? 8'hd5 : _GEN_3175; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3177 = 8'h69 == io_in_0 ? 8'hde : _GEN_3176; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3178 = 8'h6a == io_in_0 ? 8'hc3 : _GEN_3177; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3179 = 8'h6b == io_in_0 ? 8'hc8 : _GEN_3178; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3180 = 8'h6c == io_in_0 ? 8'hf9 : _GEN_3179; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3181 = 8'h6d == io_in_0 ? 8'hf2 : _GEN_3180; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3182 = 8'h6e == io_in_0 ? 8'hef : _GEN_3181; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3183 = 8'h6f == io_in_0 ? 8'he4 : _GEN_3182; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3184 = 8'h70 == io_in_0 ? 8'h3d : _GEN_3183; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3185 = 8'h71 == io_in_0 ? 8'h36 : _GEN_3184; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3186 = 8'h72 == io_in_0 ? 8'h2b : _GEN_3185; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3187 = 8'h73 == io_in_0 ? 8'h20 : _GEN_3186; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3188 = 8'h74 == io_in_0 ? 8'h11 : _GEN_3187; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3189 = 8'h75 == io_in_0 ? 8'h1a : _GEN_3188; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3190 = 8'h76 == io_in_0 ? 8'h7 : _GEN_3189; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3191 = 8'h77 == io_in_0 ? 8'hc : _GEN_3190; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3192 = 8'h78 == io_in_0 ? 8'h65 : _GEN_3191; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3193 = 8'h79 == io_in_0 ? 8'h6e : _GEN_3192; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3194 = 8'h7a == io_in_0 ? 8'h73 : _GEN_3193; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3195 = 8'h7b == io_in_0 ? 8'h78 : _GEN_3194; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3196 = 8'h7c == io_in_0 ? 8'h49 : _GEN_3195; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3197 = 8'h7d == io_in_0 ? 8'h42 : _GEN_3196; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3198 = 8'h7e == io_in_0 ? 8'h5f : _GEN_3197; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3199 = 8'h7f == io_in_0 ? 8'h54 : _GEN_3198; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3200 = 8'h80 == io_in_0 ? 8'hf7 : _GEN_3199; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3201 = 8'h81 == io_in_0 ? 8'hfc : _GEN_3200; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3202 = 8'h82 == io_in_0 ? 8'he1 : _GEN_3201; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3203 = 8'h83 == io_in_0 ? 8'hea : _GEN_3202; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3204 = 8'h84 == io_in_0 ? 8'hdb : _GEN_3203; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3205 = 8'h85 == io_in_0 ? 8'hd0 : _GEN_3204; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3206 = 8'h86 == io_in_0 ? 8'hcd : _GEN_3205; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3207 = 8'h87 == io_in_0 ? 8'hc6 : _GEN_3206; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3208 = 8'h88 == io_in_0 ? 8'haf : _GEN_3207; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3209 = 8'h89 == io_in_0 ? 8'ha4 : _GEN_3208; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3210 = 8'h8a == io_in_0 ? 8'hb9 : _GEN_3209; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3211 = 8'h8b == io_in_0 ? 8'hb2 : _GEN_3210; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3212 = 8'h8c == io_in_0 ? 8'h83 : _GEN_3211; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3213 = 8'h8d == io_in_0 ? 8'h88 : _GEN_3212; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3214 = 8'h8e == io_in_0 ? 8'h95 : _GEN_3213; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3215 = 8'h8f == io_in_0 ? 8'h9e : _GEN_3214; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3216 = 8'h90 == io_in_0 ? 8'h47 : _GEN_3215; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3217 = 8'h91 == io_in_0 ? 8'h4c : _GEN_3216; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3218 = 8'h92 == io_in_0 ? 8'h51 : _GEN_3217; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3219 = 8'h93 == io_in_0 ? 8'h5a : _GEN_3218; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3220 = 8'h94 == io_in_0 ? 8'h6b : _GEN_3219; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3221 = 8'h95 == io_in_0 ? 8'h60 : _GEN_3220; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3222 = 8'h96 == io_in_0 ? 8'h7d : _GEN_3221; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3223 = 8'h97 == io_in_0 ? 8'h76 : _GEN_3222; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3224 = 8'h98 == io_in_0 ? 8'h1f : _GEN_3223; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3225 = 8'h99 == io_in_0 ? 8'h14 : _GEN_3224; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3226 = 8'h9a == io_in_0 ? 8'h9 : _GEN_3225; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3227 = 8'h9b == io_in_0 ? 8'h2 : _GEN_3226; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3228 = 8'h9c == io_in_0 ? 8'h33 : _GEN_3227; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3229 = 8'h9d == io_in_0 ? 8'h38 : _GEN_3228; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3230 = 8'h9e == io_in_0 ? 8'h25 : _GEN_3229; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3231 = 8'h9f == io_in_0 ? 8'h2e : _GEN_3230; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3232 = 8'ha0 == io_in_0 ? 8'h8c : _GEN_3231; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3233 = 8'ha1 == io_in_0 ? 8'h87 : _GEN_3232; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3234 = 8'ha2 == io_in_0 ? 8'h9a : _GEN_3233; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3235 = 8'ha3 == io_in_0 ? 8'h91 : _GEN_3234; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3236 = 8'ha4 == io_in_0 ? 8'ha0 : _GEN_3235; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3237 = 8'ha5 == io_in_0 ? 8'hab : _GEN_3236; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3238 = 8'ha6 == io_in_0 ? 8'hb6 : _GEN_3237; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3239 = 8'ha7 == io_in_0 ? 8'hbd : _GEN_3238; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3240 = 8'ha8 == io_in_0 ? 8'hd4 : _GEN_3239; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3241 = 8'ha9 == io_in_0 ? 8'hdf : _GEN_3240; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3242 = 8'haa == io_in_0 ? 8'hc2 : _GEN_3241; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3243 = 8'hab == io_in_0 ? 8'hc9 : _GEN_3242; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3244 = 8'hac == io_in_0 ? 8'hf8 : _GEN_3243; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3245 = 8'had == io_in_0 ? 8'hf3 : _GEN_3244; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3246 = 8'hae == io_in_0 ? 8'hee : _GEN_3245; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3247 = 8'haf == io_in_0 ? 8'he5 : _GEN_3246; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3248 = 8'hb0 == io_in_0 ? 8'h3c : _GEN_3247; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3249 = 8'hb1 == io_in_0 ? 8'h37 : _GEN_3248; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3250 = 8'hb2 == io_in_0 ? 8'h2a : _GEN_3249; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3251 = 8'hb3 == io_in_0 ? 8'h21 : _GEN_3250; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3252 = 8'hb4 == io_in_0 ? 8'h10 : _GEN_3251; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3253 = 8'hb5 == io_in_0 ? 8'h1b : _GEN_3252; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3254 = 8'hb6 == io_in_0 ? 8'h6 : _GEN_3253; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3255 = 8'hb7 == io_in_0 ? 8'hd : _GEN_3254; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3256 = 8'hb8 == io_in_0 ? 8'h64 : _GEN_3255; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3257 = 8'hb9 == io_in_0 ? 8'h6f : _GEN_3256; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3258 = 8'hba == io_in_0 ? 8'h72 : _GEN_3257; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3259 = 8'hbb == io_in_0 ? 8'h79 : _GEN_3258; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3260 = 8'hbc == io_in_0 ? 8'h48 : _GEN_3259; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3261 = 8'hbd == io_in_0 ? 8'h43 : _GEN_3260; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3262 = 8'hbe == io_in_0 ? 8'h5e : _GEN_3261; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3263 = 8'hbf == io_in_0 ? 8'h55 : _GEN_3262; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3264 = 8'hc0 == io_in_0 ? 8'h1 : _GEN_3263; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3265 = 8'hc1 == io_in_0 ? 8'ha : _GEN_3264; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3266 = 8'hc2 == io_in_0 ? 8'h17 : _GEN_3265; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3267 = 8'hc3 == io_in_0 ? 8'h1c : _GEN_3266; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3268 = 8'hc4 == io_in_0 ? 8'h2d : _GEN_3267; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3269 = 8'hc5 == io_in_0 ? 8'h26 : _GEN_3268; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3270 = 8'hc6 == io_in_0 ? 8'h3b : _GEN_3269; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3271 = 8'hc7 == io_in_0 ? 8'h30 : _GEN_3270; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3272 = 8'hc8 == io_in_0 ? 8'h59 : _GEN_3271; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3273 = 8'hc9 == io_in_0 ? 8'h52 : _GEN_3272; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3274 = 8'hca == io_in_0 ? 8'h4f : _GEN_3273; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3275 = 8'hcb == io_in_0 ? 8'h44 : _GEN_3274; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3276 = 8'hcc == io_in_0 ? 8'h75 : _GEN_3275; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3277 = 8'hcd == io_in_0 ? 8'h7e : _GEN_3276; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3278 = 8'hce == io_in_0 ? 8'h63 : _GEN_3277; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3279 = 8'hcf == io_in_0 ? 8'h68 : _GEN_3278; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3280 = 8'hd0 == io_in_0 ? 8'hb1 : _GEN_3279; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3281 = 8'hd1 == io_in_0 ? 8'hba : _GEN_3280; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3282 = 8'hd2 == io_in_0 ? 8'ha7 : _GEN_3281; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3283 = 8'hd3 == io_in_0 ? 8'hac : _GEN_3282; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3284 = 8'hd4 == io_in_0 ? 8'h9d : _GEN_3283; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3285 = 8'hd5 == io_in_0 ? 8'h96 : _GEN_3284; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3286 = 8'hd6 == io_in_0 ? 8'h8b : _GEN_3285; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3287 = 8'hd7 == io_in_0 ? 8'h80 : _GEN_3286; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3288 = 8'hd8 == io_in_0 ? 8'he9 : _GEN_3287; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3289 = 8'hd9 == io_in_0 ? 8'he2 : _GEN_3288; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3290 = 8'hda == io_in_0 ? 8'hff : _GEN_3289; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3291 = 8'hdb == io_in_0 ? 8'hf4 : _GEN_3290; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3292 = 8'hdc == io_in_0 ? 8'hc5 : _GEN_3291; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3293 = 8'hdd == io_in_0 ? 8'hce : _GEN_3292; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3294 = 8'hde == io_in_0 ? 8'hd3 : _GEN_3293; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3295 = 8'hdf == io_in_0 ? 8'hd8 : _GEN_3294; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3296 = 8'he0 == io_in_0 ? 8'h7a : _GEN_3295; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3297 = 8'he1 == io_in_0 ? 8'h71 : _GEN_3296; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3298 = 8'he2 == io_in_0 ? 8'h6c : _GEN_3297; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3299 = 8'he3 == io_in_0 ? 8'h67 : _GEN_3298; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3300 = 8'he4 == io_in_0 ? 8'h56 : _GEN_3299; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3301 = 8'he5 == io_in_0 ? 8'h5d : _GEN_3300; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3302 = 8'he6 == io_in_0 ? 8'h40 : _GEN_3301; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3303 = 8'he7 == io_in_0 ? 8'h4b : _GEN_3302; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3304 = 8'he8 == io_in_0 ? 8'h22 : _GEN_3303; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3305 = 8'he9 == io_in_0 ? 8'h29 : _GEN_3304; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3306 = 8'hea == io_in_0 ? 8'h34 : _GEN_3305; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3307 = 8'heb == io_in_0 ? 8'h3f : _GEN_3306; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3308 = 8'hec == io_in_0 ? 8'he : _GEN_3307; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3309 = 8'hed == io_in_0 ? 8'h5 : _GEN_3308; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3310 = 8'hee == io_in_0 ? 8'h18 : _GEN_3309; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3311 = 8'hef == io_in_0 ? 8'h13 : _GEN_3310; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3312 = 8'hf0 == io_in_0 ? 8'hca : _GEN_3311; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3313 = 8'hf1 == io_in_0 ? 8'hc1 : _GEN_3312; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3314 = 8'hf2 == io_in_0 ? 8'hdc : _GEN_3313; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3315 = 8'hf3 == io_in_0 ? 8'hd7 : _GEN_3314; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3316 = 8'hf4 == io_in_0 ? 8'he6 : _GEN_3315; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3317 = 8'hf5 == io_in_0 ? 8'hed : _GEN_3316; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3318 = 8'hf6 == io_in_0 ? 8'hf0 : _GEN_3317; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3319 = 8'hf7 == io_in_0 ? 8'hfb : _GEN_3318; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3320 = 8'hf8 == io_in_0 ? 8'h92 : _GEN_3319; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3321 = 8'hf9 == io_in_0 ? 8'h99 : _GEN_3320; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3322 = 8'hfa == io_in_0 ? 8'h84 : _GEN_3321; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3323 = 8'hfb == io_in_0 ? 8'h8f : _GEN_3322; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3324 = 8'hfc == io_in_0 ? 8'hbe : _GEN_3323; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3325 = 8'hfd == io_in_0 ? 8'hb5 : _GEN_3324; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3326 = 8'hfe == io_in_0 ? 8'ha8 : _GEN_3325; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3327 = 8'hff == io_in_0 ? 8'ha3 : _GEN_3326; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3329 = 8'h1 == io_in_1 ? 8'hd : 8'h0; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3330 = 8'h2 == io_in_1 ? 8'h1a : _GEN_3329; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3331 = 8'h3 == io_in_1 ? 8'h17 : _GEN_3330; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3332 = 8'h4 == io_in_1 ? 8'h34 : _GEN_3331; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3333 = 8'h5 == io_in_1 ? 8'h39 : _GEN_3332; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3334 = 8'h6 == io_in_1 ? 8'h2e : _GEN_3333; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3335 = 8'h7 == io_in_1 ? 8'h23 : _GEN_3334; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3336 = 8'h8 == io_in_1 ? 8'h68 : _GEN_3335; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3337 = 8'h9 == io_in_1 ? 8'h65 : _GEN_3336; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3338 = 8'ha == io_in_1 ? 8'h72 : _GEN_3337; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3339 = 8'hb == io_in_1 ? 8'h7f : _GEN_3338; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3340 = 8'hc == io_in_1 ? 8'h5c : _GEN_3339; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3341 = 8'hd == io_in_1 ? 8'h51 : _GEN_3340; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3342 = 8'he == io_in_1 ? 8'h46 : _GEN_3341; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3343 = 8'hf == io_in_1 ? 8'h4b : _GEN_3342; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3344 = 8'h10 == io_in_1 ? 8'hd0 : _GEN_3343; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3345 = 8'h11 == io_in_1 ? 8'hdd : _GEN_3344; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3346 = 8'h12 == io_in_1 ? 8'hca : _GEN_3345; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3347 = 8'h13 == io_in_1 ? 8'hc7 : _GEN_3346; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3348 = 8'h14 == io_in_1 ? 8'he4 : _GEN_3347; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3349 = 8'h15 == io_in_1 ? 8'he9 : _GEN_3348; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3350 = 8'h16 == io_in_1 ? 8'hfe : _GEN_3349; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3351 = 8'h17 == io_in_1 ? 8'hf3 : _GEN_3350; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3352 = 8'h18 == io_in_1 ? 8'hb8 : _GEN_3351; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3353 = 8'h19 == io_in_1 ? 8'hb5 : _GEN_3352; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3354 = 8'h1a == io_in_1 ? 8'ha2 : _GEN_3353; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3355 = 8'h1b == io_in_1 ? 8'haf : _GEN_3354; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3356 = 8'h1c == io_in_1 ? 8'h8c : _GEN_3355; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3357 = 8'h1d == io_in_1 ? 8'h81 : _GEN_3356; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3358 = 8'h1e == io_in_1 ? 8'h96 : _GEN_3357; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3359 = 8'h1f == io_in_1 ? 8'h9b : _GEN_3358; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3360 = 8'h20 == io_in_1 ? 8'hbb : _GEN_3359; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3361 = 8'h21 == io_in_1 ? 8'hb6 : _GEN_3360; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3362 = 8'h22 == io_in_1 ? 8'ha1 : _GEN_3361; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3363 = 8'h23 == io_in_1 ? 8'hac : _GEN_3362; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3364 = 8'h24 == io_in_1 ? 8'h8f : _GEN_3363; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3365 = 8'h25 == io_in_1 ? 8'h82 : _GEN_3364; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3366 = 8'h26 == io_in_1 ? 8'h95 : _GEN_3365; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3367 = 8'h27 == io_in_1 ? 8'h98 : _GEN_3366; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3368 = 8'h28 == io_in_1 ? 8'hd3 : _GEN_3367; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3369 = 8'h29 == io_in_1 ? 8'hde : _GEN_3368; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3370 = 8'h2a == io_in_1 ? 8'hc9 : _GEN_3369; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3371 = 8'h2b == io_in_1 ? 8'hc4 : _GEN_3370; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3372 = 8'h2c == io_in_1 ? 8'he7 : _GEN_3371; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3373 = 8'h2d == io_in_1 ? 8'hea : _GEN_3372; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3374 = 8'h2e == io_in_1 ? 8'hfd : _GEN_3373; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3375 = 8'h2f == io_in_1 ? 8'hf0 : _GEN_3374; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3376 = 8'h30 == io_in_1 ? 8'h6b : _GEN_3375; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3377 = 8'h31 == io_in_1 ? 8'h66 : _GEN_3376; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3378 = 8'h32 == io_in_1 ? 8'h71 : _GEN_3377; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3379 = 8'h33 == io_in_1 ? 8'h7c : _GEN_3378; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3380 = 8'h34 == io_in_1 ? 8'h5f : _GEN_3379; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3381 = 8'h35 == io_in_1 ? 8'h52 : _GEN_3380; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3382 = 8'h36 == io_in_1 ? 8'h45 : _GEN_3381; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3383 = 8'h37 == io_in_1 ? 8'h48 : _GEN_3382; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3384 = 8'h38 == io_in_1 ? 8'h3 : _GEN_3383; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3385 = 8'h39 == io_in_1 ? 8'he : _GEN_3384; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3386 = 8'h3a == io_in_1 ? 8'h19 : _GEN_3385; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3387 = 8'h3b == io_in_1 ? 8'h14 : _GEN_3386; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3388 = 8'h3c == io_in_1 ? 8'h37 : _GEN_3387; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3389 = 8'h3d == io_in_1 ? 8'h3a : _GEN_3388; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3390 = 8'h3e == io_in_1 ? 8'h2d : _GEN_3389; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3391 = 8'h3f == io_in_1 ? 8'h20 : _GEN_3390; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3392 = 8'h40 == io_in_1 ? 8'h6d : _GEN_3391; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3393 = 8'h41 == io_in_1 ? 8'h60 : _GEN_3392; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3394 = 8'h42 == io_in_1 ? 8'h77 : _GEN_3393; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3395 = 8'h43 == io_in_1 ? 8'h7a : _GEN_3394; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3396 = 8'h44 == io_in_1 ? 8'h59 : _GEN_3395; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3397 = 8'h45 == io_in_1 ? 8'h54 : _GEN_3396; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3398 = 8'h46 == io_in_1 ? 8'h43 : _GEN_3397; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3399 = 8'h47 == io_in_1 ? 8'h4e : _GEN_3398; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3400 = 8'h48 == io_in_1 ? 8'h5 : _GEN_3399; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3401 = 8'h49 == io_in_1 ? 8'h8 : _GEN_3400; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3402 = 8'h4a == io_in_1 ? 8'h1f : _GEN_3401; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3403 = 8'h4b == io_in_1 ? 8'h12 : _GEN_3402; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3404 = 8'h4c == io_in_1 ? 8'h31 : _GEN_3403; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3405 = 8'h4d == io_in_1 ? 8'h3c : _GEN_3404; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3406 = 8'h4e == io_in_1 ? 8'h2b : _GEN_3405; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3407 = 8'h4f == io_in_1 ? 8'h26 : _GEN_3406; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3408 = 8'h50 == io_in_1 ? 8'hbd : _GEN_3407; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3409 = 8'h51 == io_in_1 ? 8'hb0 : _GEN_3408; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3410 = 8'h52 == io_in_1 ? 8'ha7 : _GEN_3409; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3411 = 8'h53 == io_in_1 ? 8'haa : _GEN_3410; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3412 = 8'h54 == io_in_1 ? 8'h89 : _GEN_3411; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3413 = 8'h55 == io_in_1 ? 8'h84 : _GEN_3412; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3414 = 8'h56 == io_in_1 ? 8'h93 : _GEN_3413; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3415 = 8'h57 == io_in_1 ? 8'h9e : _GEN_3414; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3416 = 8'h58 == io_in_1 ? 8'hd5 : _GEN_3415; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3417 = 8'h59 == io_in_1 ? 8'hd8 : _GEN_3416; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3418 = 8'h5a == io_in_1 ? 8'hcf : _GEN_3417; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3419 = 8'h5b == io_in_1 ? 8'hc2 : _GEN_3418; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3420 = 8'h5c == io_in_1 ? 8'he1 : _GEN_3419; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3421 = 8'h5d == io_in_1 ? 8'hec : _GEN_3420; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3422 = 8'h5e == io_in_1 ? 8'hfb : _GEN_3421; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3423 = 8'h5f == io_in_1 ? 8'hf6 : _GEN_3422; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3424 = 8'h60 == io_in_1 ? 8'hd6 : _GEN_3423; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3425 = 8'h61 == io_in_1 ? 8'hdb : _GEN_3424; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3426 = 8'h62 == io_in_1 ? 8'hcc : _GEN_3425; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3427 = 8'h63 == io_in_1 ? 8'hc1 : _GEN_3426; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3428 = 8'h64 == io_in_1 ? 8'he2 : _GEN_3427; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3429 = 8'h65 == io_in_1 ? 8'hef : _GEN_3428; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3430 = 8'h66 == io_in_1 ? 8'hf8 : _GEN_3429; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3431 = 8'h67 == io_in_1 ? 8'hf5 : _GEN_3430; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3432 = 8'h68 == io_in_1 ? 8'hbe : _GEN_3431; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3433 = 8'h69 == io_in_1 ? 8'hb3 : _GEN_3432; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3434 = 8'h6a == io_in_1 ? 8'ha4 : _GEN_3433; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3435 = 8'h6b == io_in_1 ? 8'ha9 : _GEN_3434; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3436 = 8'h6c == io_in_1 ? 8'h8a : _GEN_3435; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3437 = 8'h6d == io_in_1 ? 8'h87 : _GEN_3436; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3438 = 8'h6e == io_in_1 ? 8'h90 : _GEN_3437; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3439 = 8'h6f == io_in_1 ? 8'h9d : _GEN_3438; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3440 = 8'h70 == io_in_1 ? 8'h6 : _GEN_3439; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3441 = 8'h71 == io_in_1 ? 8'hb : _GEN_3440; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3442 = 8'h72 == io_in_1 ? 8'h1c : _GEN_3441; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3443 = 8'h73 == io_in_1 ? 8'h11 : _GEN_3442; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3444 = 8'h74 == io_in_1 ? 8'h32 : _GEN_3443; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3445 = 8'h75 == io_in_1 ? 8'h3f : _GEN_3444; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3446 = 8'h76 == io_in_1 ? 8'h28 : _GEN_3445; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3447 = 8'h77 == io_in_1 ? 8'h25 : _GEN_3446; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3448 = 8'h78 == io_in_1 ? 8'h6e : _GEN_3447; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3449 = 8'h79 == io_in_1 ? 8'h63 : _GEN_3448; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3450 = 8'h7a == io_in_1 ? 8'h74 : _GEN_3449; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3451 = 8'h7b == io_in_1 ? 8'h79 : _GEN_3450; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3452 = 8'h7c == io_in_1 ? 8'h5a : _GEN_3451; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3453 = 8'h7d == io_in_1 ? 8'h57 : _GEN_3452; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3454 = 8'h7e == io_in_1 ? 8'h40 : _GEN_3453; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3455 = 8'h7f == io_in_1 ? 8'h4d : _GEN_3454; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3456 = 8'h80 == io_in_1 ? 8'hda : _GEN_3455; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3457 = 8'h81 == io_in_1 ? 8'hd7 : _GEN_3456; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3458 = 8'h82 == io_in_1 ? 8'hc0 : _GEN_3457; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3459 = 8'h83 == io_in_1 ? 8'hcd : _GEN_3458; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3460 = 8'h84 == io_in_1 ? 8'hee : _GEN_3459; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3461 = 8'h85 == io_in_1 ? 8'he3 : _GEN_3460; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3462 = 8'h86 == io_in_1 ? 8'hf4 : _GEN_3461; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3463 = 8'h87 == io_in_1 ? 8'hf9 : _GEN_3462; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3464 = 8'h88 == io_in_1 ? 8'hb2 : _GEN_3463; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3465 = 8'h89 == io_in_1 ? 8'hbf : _GEN_3464; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3466 = 8'h8a == io_in_1 ? 8'ha8 : _GEN_3465; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3467 = 8'h8b == io_in_1 ? 8'ha5 : _GEN_3466; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3468 = 8'h8c == io_in_1 ? 8'h86 : _GEN_3467; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3469 = 8'h8d == io_in_1 ? 8'h8b : _GEN_3468; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3470 = 8'h8e == io_in_1 ? 8'h9c : _GEN_3469; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3471 = 8'h8f == io_in_1 ? 8'h91 : _GEN_3470; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3472 = 8'h90 == io_in_1 ? 8'ha : _GEN_3471; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3473 = 8'h91 == io_in_1 ? 8'h7 : _GEN_3472; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3474 = 8'h92 == io_in_1 ? 8'h10 : _GEN_3473; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3475 = 8'h93 == io_in_1 ? 8'h1d : _GEN_3474; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3476 = 8'h94 == io_in_1 ? 8'h3e : _GEN_3475; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3477 = 8'h95 == io_in_1 ? 8'h33 : _GEN_3476; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3478 = 8'h96 == io_in_1 ? 8'h24 : _GEN_3477; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3479 = 8'h97 == io_in_1 ? 8'h29 : _GEN_3478; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3480 = 8'h98 == io_in_1 ? 8'h62 : _GEN_3479; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3481 = 8'h99 == io_in_1 ? 8'h6f : _GEN_3480; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3482 = 8'h9a == io_in_1 ? 8'h78 : _GEN_3481; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3483 = 8'h9b == io_in_1 ? 8'h75 : _GEN_3482; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3484 = 8'h9c == io_in_1 ? 8'h56 : _GEN_3483; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3485 = 8'h9d == io_in_1 ? 8'h5b : _GEN_3484; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3486 = 8'h9e == io_in_1 ? 8'h4c : _GEN_3485; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3487 = 8'h9f == io_in_1 ? 8'h41 : _GEN_3486; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3488 = 8'ha0 == io_in_1 ? 8'h61 : _GEN_3487; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3489 = 8'ha1 == io_in_1 ? 8'h6c : _GEN_3488; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3490 = 8'ha2 == io_in_1 ? 8'h7b : _GEN_3489; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3491 = 8'ha3 == io_in_1 ? 8'h76 : _GEN_3490; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3492 = 8'ha4 == io_in_1 ? 8'h55 : _GEN_3491; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3493 = 8'ha5 == io_in_1 ? 8'h58 : _GEN_3492; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3494 = 8'ha6 == io_in_1 ? 8'h4f : _GEN_3493; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3495 = 8'ha7 == io_in_1 ? 8'h42 : _GEN_3494; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3496 = 8'ha8 == io_in_1 ? 8'h9 : _GEN_3495; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3497 = 8'ha9 == io_in_1 ? 8'h4 : _GEN_3496; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3498 = 8'haa == io_in_1 ? 8'h13 : _GEN_3497; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3499 = 8'hab == io_in_1 ? 8'h1e : _GEN_3498; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3500 = 8'hac == io_in_1 ? 8'h3d : _GEN_3499; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3501 = 8'had == io_in_1 ? 8'h30 : _GEN_3500; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3502 = 8'hae == io_in_1 ? 8'h27 : _GEN_3501; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3503 = 8'haf == io_in_1 ? 8'h2a : _GEN_3502; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3504 = 8'hb0 == io_in_1 ? 8'hb1 : _GEN_3503; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3505 = 8'hb1 == io_in_1 ? 8'hbc : _GEN_3504; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3506 = 8'hb2 == io_in_1 ? 8'hab : _GEN_3505; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3507 = 8'hb3 == io_in_1 ? 8'ha6 : _GEN_3506; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3508 = 8'hb4 == io_in_1 ? 8'h85 : _GEN_3507; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3509 = 8'hb5 == io_in_1 ? 8'h88 : _GEN_3508; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3510 = 8'hb6 == io_in_1 ? 8'h9f : _GEN_3509; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3511 = 8'hb7 == io_in_1 ? 8'h92 : _GEN_3510; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3512 = 8'hb8 == io_in_1 ? 8'hd9 : _GEN_3511; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3513 = 8'hb9 == io_in_1 ? 8'hd4 : _GEN_3512; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3514 = 8'hba == io_in_1 ? 8'hc3 : _GEN_3513; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3515 = 8'hbb == io_in_1 ? 8'hce : _GEN_3514; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3516 = 8'hbc == io_in_1 ? 8'hed : _GEN_3515; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3517 = 8'hbd == io_in_1 ? 8'he0 : _GEN_3516; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3518 = 8'hbe == io_in_1 ? 8'hf7 : _GEN_3517; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3519 = 8'hbf == io_in_1 ? 8'hfa : _GEN_3518; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3520 = 8'hc0 == io_in_1 ? 8'hb7 : _GEN_3519; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3521 = 8'hc1 == io_in_1 ? 8'hba : _GEN_3520; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3522 = 8'hc2 == io_in_1 ? 8'had : _GEN_3521; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3523 = 8'hc3 == io_in_1 ? 8'ha0 : _GEN_3522; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3524 = 8'hc4 == io_in_1 ? 8'h83 : _GEN_3523; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3525 = 8'hc5 == io_in_1 ? 8'h8e : _GEN_3524; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3526 = 8'hc6 == io_in_1 ? 8'h99 : _GEN_3525; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3527 = 8'hc7 == io_in_1 ? 8'h94 : _GEN_3526; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3528 = 8'hc8 == io_in_1 ? 8'hdf : _GEN_3527; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3529 = 8'hc9 == io_in_1 ? 8'hd2 : _GEN_3528; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3530 = 8'hca == io_in_1 ? 8'hc5 : _GEN_3529; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3531 = 8'hcb == io_in_1 ? 8'hc8 : _GEN_3530; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3532 = 8'hcc == io_in_1 ? 8'heb : _GEN_3531; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3533 = 8'hcd == io_in_1 ? 8'he6 : _GEN_3532; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3534 = 8'hce == io_in_1 ? 8'hf1 : _GEN_3533; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3535 = 8'hcf == io_in_1 ? 8'hfc : _GEN_3534; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3536 = 8'hd0 == io_in_1 ? 8'h67 : _GEN_3535; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3537 = 8'hd1 == io_in_1 ? 8'h6a : _GEN_3536; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3538 = 8'hd2 == io_in_1 ? 8'h7d : _GEN_3537; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3539 = 8'hd3 == io_in_1 ? 8'h70 : _GEN_3538; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3540 = 8'hd4 == io_in_1 ? 8'h53 : _GEN_3539; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3541 = 8'hd5 == io_in_1 ? 8'h5e : _GEN_3540; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3542 = 8'hd6 == io_in_1 ? 8'h49 : _GEN_3541; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3543 = 8'hd7 == io_in_1 ? 8'h44 : _GEN_3542; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3544 = 8'hd8 == io_in_1 ? 8'hf : _GEN_3543; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3545 = 8'hd9 == io_in_1 ? 8'h2 : _GEN_3544; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3546 = 8'hda == io_in_1 ? 8'h15 : _GEN_3545; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3547 = 8'hdb == io_in_1 ? 8'h18 : _GEN_3546; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3548 = 8'hdc == io_in_1 ? 8'h3b : _GEN_3547; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3549 = 8'hdd == io_in_1 ? 8'h36 : _GEN_3548; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3550 = 8'hde == io_in_1 ? 8'h21 : _GEN_3549; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3551 = 8'hdf == io_in_1 ? 8'h2c : _GEN_3550; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3552 = 8'he0 == io_in_1 ? 8'hc : _GEN_3551; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3553 = 8'he1 == io_in_1 ? 8'h1 : _GEN_3552; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3554 = 8'he2 == io_in_1 ? 8'h16 : _GEN_3553; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3555 = 8'he3 == io_in_1 ? 8'h1b : _GEN_3554; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3556 = 8'he4 == io_in_1 ? 8'h38 : _GEN_3555; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3557 = 8'he5 == io_in_1 ? 8'h35 : _GEN_3556; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3558 = 8'he6 == io_in_1 ? 8'h22 : _GEN_3557; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3559 = 8'he7 == io_in_1 ? 8'h2f : _GEN_3558; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3560 = 8'he8 == io_in_1 ? 8'h64 : _GEN_3559; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3561 = 8'he9 == io_in_1 ? 8'h69 : _GEN_3560; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3562 = 8'hea == io_in_1 ? 8'h7e : _GEN_3561; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3563 = 8'heb == io_in_1 ? 8'h73 : _GEN_3562; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3564 = 8'hec == io_in_1 ? 8'h50 : _GEN_3563; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3565 = 8'hed == io_in_1 ? 8'h5d : _GEN_3564; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3566 = 8'hee == io_in_1 ? 8'h4a : _GEN_3565; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3567 = 8'hef == io_in_1 ? 8'h47 : _GEN_3566; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3568 = 8'hf0 == io_in_1 ? 8'hdc : _GEN_3567; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3569 = 8'hf1 == io_in_1 ? 8'hd1 : _GEN_3568; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3570 = 8'hf2 == io_in_1 ? 8'hc6 : _GEN_3569; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3571 = 8'hf3 == io_in_1 ? 8'hcb : _GEN_3570; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3572 = 8'hf4 == io_in_1 ? 8'he8 : _GEN_3571; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3573 = 8'hf5 == io_in_1 ? 8'he5 : _GEN_3572; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3574 = 8'hf6 == io_in_1 ? 8'hf2 : _GEN_3573; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3575 = 8'hf7 == io_in_1 ? 8'hff : _GEN_3574; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3576 = 8'hf8 == io_in_1 ? 8'hb4 : _GEN_3575; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3577 = 8'hf9 == io_in_1 ? 8'hb9 : _GEN_3576; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3578 = 8'hfa == io_in_1 ? 8'hae : _GEN_3577; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3579 = 8'hfb == io_in_1 ? 8'ha3 : _GEN_3578; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3580 = 8'hfc == io_in_1 ? 8'h80 : _GEN_3579; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3581 = 8'hfd == io_in_1 ? 8'h8d : _GEN_3580; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3582 = 8'hfe == io_in_1 ? 8'h9a : _GEN_3581; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3583 = 8'hff == io_in_1 ? 8'h97 : _GEN_3582; // @[AES_PipelinedElasticBuffer.scala 594:32 AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _T_9 = _GEN_3327 ^ _GEN_3583; // @[AES_PipelinedElasticBuffer.scala 594:32]
  wire [7:0] _GEN_3585 = 8'h1 == io_in_2 ? 8'h9 : 8'h0; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3586 = 8'h2 == io_in_2 ? 8'h12 : _GEN_3585; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3587 = 8'h3 == io_in_2 ? 8'h1b : _GEN_3586; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3588 = 8'h4 == io_in_2 ? 8'h24 : _GEN_3587; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3589 = 8'h5 == io_in_2 ? 8'h2d : _GEN_3588; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3590 = 8'h6 == io_in_2 ? 8'h36 : _GEN_3589; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3591 = 8'h7 == io_in_2 ? 8'h3f : _GEN_3590; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3592 = 8'h8 == io_in_2 ? 8'h48 : _GEN_3591; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3593 = 8'h9 == io_in_2 ? 8'h41 : _GEN_3592; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3594 = 8'ha == io_in_2 ? 8'h5a : _GEN_3593; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3595 = 8'hb == io_in_2 ? 8'h53 : _GEN_3594; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3596 = 8'hc == io_in_2 ? 8'h6c : _GEN_3595; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3597 = 8'hd == io_in_2 ? 8'h65 : _GEN_3596; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3598 = 8'he == io_in_2 ? 8'h7e : _GEN_3597; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3599 = 8'hf == io_in_2 ? 8'h77 : _GEN_3598; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3600 = 8'h10 == io_in_2 ? 8'h90 : _GEN_3599; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3601 = 8'h11 == io_in_2 ? 8'h99 : _GEN_3600; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3602 = 8'h12 == io_in_2 ? 8'h82 : _GEN_3601; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3603 = 8'h13 == io_in_2 ? 8'h8b : _GEN_3602; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3604 = 8'h14 == io_in_2 ? 8'hb4 : _GEN_3603; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3605 = 8'h15 == io_in_2 ? 8'hbd : _GEN_3604; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3606 = 8'h16 == io_in_2 ? 8'ha6 : _GEN_3605; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3607 = 8'h17 == io_in_2 ? 8'haf : _GEN_3606; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3608 = 8'h18 == io_in_2 ? 8'hd8 : _GEN_3607; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3609 = 8'h19 == io_in_2 ? 8'hd1 : _GEN_3608; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3610 = 8'h1a == io_in_2 ? 8'hca : _GEN_3609; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3611 = 8'h1b == io_in_2 ? 8'hc3 : _GEN_3610; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3612 = 8'h1c == io_in_2 ? 8'hfc : _GEN_3611; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3613 = 8'h1d == io_in_2 ? 8'hf5 : _GEN_3612; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3614 = 8'h1e == io_in_2 ? 8'hee : _GEN_3613; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3615 = 8'h1f == io_in_2 ? 8'he7 : _GEN_3614; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3616 = 8'h20 == io_in_2 ? 8'h3b : _GEN_3615; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3617 = 8'h21 == io_in_2 ? 8'h32 : _GEN_3616; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3618 = 8'h22 == io_in_2 ? 8'h29 : _GEN_3617; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3619 = 8'h23 == io_in_2 ? 8'h20 : _GEN_3618; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3620 = 8'h24 == io_in_2 ? 8'h1f : _GEN_3619; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3621 = 8'h25 == io_in_2 ? 8'h16 : _GEN_3620; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3622 = 8'h26 == io_in_2 ? 8'hd : _GEN_3621; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3623 = 8'h27 == io_in_2 ? 8'h4 : _GEN_3622; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3624 = 8'h28 == io_in_2 ? 8'h73 : _GEN_3623; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3625 = 8'h29 == io_in_2 ? 8'h7a : _GEN_3624; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3626 = 8'h2a == io_in_2 ? 8'h61 : _GEN_3625; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3627 = 8'h2b == io_in_2 ? 8'h68 : _GEN_3626; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3628 = 8'h2c == io_in_2 ? 8'h57 : _GEN_3627; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3629 = 8'h2d == io_in_2 ? 8'h5e : _GEN_3628; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3630 = 8'h2e == io_in_2 ? 8'h45 : _GEN_3629; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3631 = 8'h2f == io_in_2 ? 8'h4c : _GEN_3630; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3632 = 8'h30 == io_in_2 ? 8'hab : _GEN_3631; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3633 = 8'h31 == io_in_2 ? 8'ha2 : _GEN_3632; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3634 = 8'h32 == io_in_2 ? 8'hb9 : _GEN_3633; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3635 = 8'h33 == io_in_2 ? 8'hb0 : _GEN_3634; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3636 = 8'h34 == io_in_2 ? 8'h8f : _GEN_3635; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3637 = 8'h35 == io_in_2 ? 8'h86 : _GEN_3636; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3638 = 8'h36 == io_in_2 ? 8'h9d : _GEN_3637; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3639 = 8'h37 == io_in_2 ? 8'h94 : _GEN_3638; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3640 = 8'h38 == io_in_2 ? 8'he3 : _GEN_3639; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3641 = 8'h39 == io_in_2 ? 8'hea : _GEN_3640; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3642 = 8'h3a == io_in_2 ? 8'hf1 : _GEN_3641; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3643 = 8'h3b == io_in_2 ? 8'hf8 : _GEN_3642; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3644 = 8'h3c == io_in_2 ? 8'hc7 : _GEN_3643; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3645 = 8'h3d == io_in_2 ? 8'hce : _GEN_3644; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3646 = 8'h3e == io_in_2 ? 8'hd5 : _GEN_3645; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3647 = 8'h3f == io_in_2 ? 8'hdc : _GEN_3646; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3648 = 8'h40 == io_in_2 ? 8'h76 : _GEN_3647; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3649 = 8'h41 == io_in_2 ? 8'h7f : _GEN_3648; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3650 = 8'h42 == io_in_2 ? 8'h64 : _GEN_3649; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3651 = 8'h43 == io_in_2 ? 8'h6d : _GEN_3650; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3652 = 8'h44 == io_in_2 ? 8'h52 : _GEN_3651; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3653 = 8'h45 == io_in_2 ? 8'h5b : _GEN_3652; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3654 = 8'h46 == io_in_2 ? 8'h40 : _GEN_3653; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3655 = 8'h47 == io_in_2 ? 8'h49 : _GEN_3654; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3656 = 8'h48 == io_in_2 ? 8'h3e : _GEN_3655; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3657 = 8'h49 == io_in_2 ? 8'h37 : _GEN_3656; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3658 = 8'h4a == io_in_2 ? 8'h2c : _GEN_3657; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3659 = 8'h4b == io_in_2 ? 8'h25 : _GEN_3658; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3660 = 8'h4c == io_in_2 ? 8'h1a : _GEN_3659; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3661 = 8'h4d == io_in_2 ? 8'h13 : _GEN_3660; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3662 = 8'h4e == io_in_2 ? 8'h8 : _GEN_3661; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3663 = 8'h4f == io_in_2 ? 8'h1 : _GEN_3662; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3664 = 8'h50 == io_in_2 ? 8'he6 : _GEN_3663; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3665 = 8'h51 == io_in_2 ? 8'hef : _GEN_3664; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3666 = 8'h52 == io_in_2 ? 8'hf4 : _GEN_3665; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3667 = 8'h53 == io_in_2 ? 8'hfd : _GEN_3666; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3668 = 8'h54 == io_in_2 ? 8'hc2 : _GEN_3667; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3669 = 8'h55 == io_in_2 ? 8'hcb : _GEN_3668; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3670 = 8'h56 == io_in_2 ? 8'hd0 : _GEN_3669; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3671 = 8'h57 == io_in_2 ? 8'hd9 : _GEN_3670; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3672 = 8'h58 == io_in_2 ? 8'hae : _GEN_3671; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3673 = 8'h59 == io_in_2 ? 8'ha7 : _GEN_3672; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3674 = 8'h5a == io_in_2 ? 8'hbc : _GEN_3673; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3675 = 8'h5b == io_in_2 ? 8'hb5 : _GEN_3674; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3676 = 8'h5c == io_in_2 ? 8'h8a : _GEN_3675; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3677 = 8'h5d == io_in_2 ? 8'h83 : _GEN_3676; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3678 = 8'h5e == io_in_2 ? 8'h98 : _GEN_3677; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3679 = 8'h5f == io_in_2 ? 8'h91 : _GEN_3678; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3680 = 8'h60 == io_in_2 ? 8'h4d : _GEN_3679; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3681 = 8'h61 == io_in_2 ? 8'h44 : _GEN_3680; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3682 = 8'h62 == io_in_2 ? 8'h5f : _GEN_3681; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3683 = 8'h63 == io_in_2 ? 8'h56 : _GEN_3682; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3684 = 8'h64 == io_in_2 ? 8'h69 : _GEN_3683; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3685 = 8'h65 == io_in_2 ? 8'h60 : _GEN_3684; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3686 = 8'h66 == io_in_2 ? 8'h7b : _GEN_3685; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3687 = 8'h67 == io_in_2 ? 8'h72 : _GEN_3686; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3688 = 8'h68 == io_in_2 ? 8'h5 : _GEN_3687; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3689 = 8'h69 == io_in_2 ? 8'hc : _GEN_3688; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3690 = 8'h6a == io_in_2 ? 8'h17 : _GEN_3689; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3691 = 8'h6b == io_in_2 ? 8'h1e : _GEN_3690; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3692 = 8'h6c == io_in_2 ? 8'h21 : _GEN_3691; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3693 = 8'h6d == io_in_2 ? 8'h28 : _GEN_3692; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3694 = 8'h6e == io_in_2 ? 8'h33 : _GEN_3693; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3695 = 8'h6f == io_in_2 ? 8'h3a : _GEN_3694; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3696 = 8'h70 == io_in_2 ? 8'hdd : _GEN_3695; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3697 = 8'h71 == io_in_2 ? 8'hd4 : _GEN_3696; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3698 = 8'h72 == io_in_2 ? 8'hcf : _GEN_3697; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3699 = 8'h73 == io_in_2 ? 8'hc6 : _GEN_3698; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3700 = 8'h74 == io_in_2 ? 8'hf9 : _GEN_3699; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3701 = 8'h75 == io_in_2 ? 8'hf0 : _GEN_3700; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3702 = 8'h76 == io_in_2 ? 8'heb : _GEN_3701; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3703 = 8'h77 == io_in_2 ? 8'he2 : _GEN_3702; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3704 = 8'h78 == io_in_2 ? 8'h95 : _GEN_3703; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3705 = 8'h79 == io_in_2 ? 8'h9c : _GEN_3704; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3706 = 8'h7a == io_in_2 ? 8'h87 : _GEN_3705; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3707 = 8'h7b == io_in_2 ? 8'h8e : _GEN_3706; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3708 = 8'h7c == io_in_2 ? 8'hb1 : _GEN_3707; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3709 = 8'h7d == io_in_2 ? 8'hb8 : _GEN_3708; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3710 = 8'h7e == io_in_2 ? 8'ha3 : _GEN_3709; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3711 = 8'h7f == io_in_2 ? 8'haa : _GEN_3710; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3712 = 8'h80 == io_in_2 ? 8'hec : _GEN_3711; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3713 = 8'h81 == io_in_2 ? 8'he5 : _GEN_3712; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3714 = 8'h82 == io_in_2 ? 8'hfe : _GEN_3713; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3715 = 8'h83 == io_in_2 ? 8'hf7 : _GEN_3714; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3716 = 8'h84 == io_in_2 ? 8'hc8 : _GEN_3715; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3717 = 8'h85 == io_in_2 ? 8'hc1 : _GEN_3716; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3718 = 8'h86 == io_in_2 ? 8'hda : _GEN_3717; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3719 = 8'h87 == io_in_2 ? 8'hd3 : _GEN_3718; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3720 = 8'h88 == io_in_2 ? 8'ha4 : _GEN_3719; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3721 = 8'h89 == io_in_2 ? 8'had : _GEN_3720; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3722 = 8'h8a == io_in_2 ? 8'hb6 : _GEN_3721; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3723 = 8'h8b == io_in_2 ? 8'hbf : _GEN_3722; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3724 = 8'h8c == io_in_2 ? 8'h80 : _GEN_3723; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3725 = 8'h8d == io_in_2 ? 8'h89 : _GEN_3724; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3726 = 8'h8e == io_in_2 ? 8'h92 : _GEN_3725; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3727 = 8'h8f == io_in_2 ? 8'h9b : _GEN_3726; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3728 = 8'h90 == io_in_2 ? 8'h7c : _GEN_3727; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3729 = 8'h91 == io_in_2 ? 8'h75 : _GEN_3728; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3730 = 8'h92 == io_in_2 ? 8'h6e : _GEN_3729; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3731 = 8'h93 == io_in_2 ? 8'h67 : _GEN_3730; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3732 = 8'h94 == io_in_2 ? 8'h58 : _GEN_3731; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3733 = 8'h95 == io_in_2 ? 8'h51 : _GEN_3732; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3734 = 8'h96 == io_in_2 ? 8'h4a : _GEN_3733; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3735 = 8'h97 == io_in_2 ? 8'h43 : _GEN_3734; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3736 = 8'h98 == io_in_2 ? 8'h34 : _GEN_3735; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3737 = 8'h99 == io_in_2 ? 8'h3d : _GEN_3736; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3738 = 8'h9a == io_in_2 ? 8'h26 : _GEN_3737; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3739 = 8'h9b == io_in_2 ? 8'h2f : _GEN_3738; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3740 = 8'h9c == io_in_2 ? 8'h10 : _GEN_3739; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3741 = 8'h9d == io_in_2 ? 8'h19 : _GEN_3740; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3742 = 8'h9e == io_in_2 ? 8'h2 : _GEN_3741; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3743 = 8'h9f == io_in_2 ? 8'hb : _GEN_3742; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3744 = 8'ha0 == io_in_2 ? 8'hd7 : _GEN_3743; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3745 = 8'ha1 == io_in_2 ? 8'hde : _GEN_3744; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3746 = 8'ha2 == io_in_2 ? 8'hc5 : _GEN_3745; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3747 = 8'ha3 == io_in_2 ? 8'hcc : _GEN_3746; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3748 = 8'ha4 == io_in_2 ? 8'hf3 : _GEN_3747; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3749 = 8'ha5 == io_in_2 ? 8'hfa : _GEN_3748; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3750 = 8'ha6 == io_in_2 ? 8'he1 : _GEN_3749; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3751 = 8'ha7 == io_in_2 ? 8'he8 : _GEN_3750; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3752 = 8'ha8 == io_in_2 ? 8'h9f : _GEN_3751; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3753 = 8'ha9 == io_in_2 ? 8'h96 : _GEN_3752; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3754 = 8'haa == io_in_2 ? 8'h8d : _GEN_3753; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3755 = 8'hab == io_in_2 ? 8'h84 : _GEN_3754; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3756 = 8'hac == io_in_2 ? 8'hbb : _GEN_3755; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3757 = 8'had == io_in_2 ? 8'hb2 : _GEN_3756; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3758 = 8'hae == io_in_2 ? 8'ha9 : _GEN_3757; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3759 = 8'haf == io_in_2 ? 8'ha0 : _GEN_3758; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3760 = 8'hb0 == io_in_2 ? 8'h47 : _GEN_3759; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3761 = 8'hb1 == io_in_2 ? 8'h4e : _GEN_3760; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3762 = 8'hb2 == io_in_2 ? 8'h55 : _GEN_3761; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3763 = 8'hb3 == io_in_2 ? 8'h5c : _GEN_3762; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3764 = 8'hb4 == io_in_2 ? 8'h63 : _GEN_3763; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3765 = 8'hb5 == io_in_2 ? 8'h6a : _GEN_3764; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3766 = 8'hb6 == io_in_2 ? 8'h71 : _GEN_3765; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3767 = 8'hb7 == io_in_2 ? 8'h78 : _GEN_3766; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3768 = 8'hb8 == io_in_2 ? 8'hf : _GEN_3767; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3769 = 8'hb9 == io_in_2 ? 8'h6 : _GEN_3768; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3770 = 8'hba == io_in_2 ? 8'h1d : _GEN_3769; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3771 = 8'hbb == io_in_2 ? 8'h14 : _GEN_3770; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3772 = 8'hbc == io_in_2 ? 8'h2b : _GEN_3771; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3773 = 8'hbd == io_in_2 ? 8'h22 : _GEN_3772; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3774 = 8'hbe == io_in_2 ? 8'h39 : _GEN_3773; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3775 = 8'hbf == io_in_2 ? 8'h30 : _GEN_3774; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3776 = 8'hc0 == io_in_2 ? 8'h9a : _GEN_3775; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3777 = 8'hc1 == io_in_2 ? 8'h93 : _GEN_3776; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3778 = 8'hc2 == io_in_2 ? 8'h88 : _GEN_3777; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3779 = 8'hc3 == io_in_2 ? 8'h81 : _GEN_3778; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3780 = 8'hc4 == io_in_2 ? 8'hbe : _GEN_3779; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3781 = 8'hc5 == io_in_2 ? 8'hb7 : _GEN_3780; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3782 = 8'hc6 == io_in_2 ? 8'hac : _GEN_3781; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3783 = 8'hc7 == io_in_2 ? 8'ha5 : _GEN_3782; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3784 = 8'hc8 == io_in_2 ? 8'hd2 : _GEN_3783; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3785 = 8'hc9 == io_in_2 ? 8'hdb : _GEN_3784; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3786 = 8'hca == io_in_2 ? 8'hc0 : _GEN_3785; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3787 = 8'hcb == io_in_2 ? 8'hc9 : _GEN_3786; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3788 = 8'hcc == io_in_2 ? 8'hf6 : _GEN_3787; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3789 = 8'hcd == io_in_2 ? 8'hff : _GEN_3788; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3790 = 8'hce == io_in_2 ? 8'he4 : _GEN_3789; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3791 = 8'hcf == io_in_2 ? 8'hed : _GEN_3790; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3792 = 8'hd0 == io_in_2 ? 8'ha : _GEN_3791; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3793 = 8'hd1 == io_in_2 ? 8'h3 : _GEN_3792; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3794 = 8'hd2 == io_in_2 ? 8'h18 : _GEN_3793; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3795 = 8'hd3 == io_in_2 ? 8'h11 : _GEN_3794; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3796 = 8'hd4 == io_in_2 ? 8'h2e : _GEN_3795; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3797 = 8'hd5 == io_in_2 ? 8'h27 : _GEN_3796; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3798 = 8'hd6 == io_in_2 ? 8'h3c : _GEN_3797; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3799 = 8'hd7 == io_in_2 ? 8'h35 : _GEN_3798; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3800 = 8'hd8 == io_in_2 ? 8'h42 : _GEN_3799; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3801 = 8'hd9 == io_in_2 ? 8'h4b : _GEN_3800; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3802 = 8'hda == io_in_2 ? 8'h50 : _GEN_3801; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3803 = 8'hdb == io_in_2 ? 8'h59 : _GEN_3802; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3804 = 8'hdc == io_in_2 ? 8'h66 : _GEN_3803; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3805 = 8'hdd == io_in_2 ? 8'h6f : _GEN_3804; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3806 = 8'hde == io_in_2 ? 8'h74 : _GEN_3805; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3807 = 8'hdf == io_in_2 ? 8'h7d : _GEN_3806; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3808 = 8'he0 == io_in_2 ? 8'ha1 : _GEN_3807; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3809 = 8'he1 == io_in_2 ? 8'ha8 : _GEN_3808; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3810 = 8'he2 == io_in_2 ? 8'hb3 : _GEN_3809; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3811 = 8'he3 == io_in_2 ? 8'hba : _GEN_3810; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3812 = 8'he4 == io_in_2 ? 8'h85 : _GEN_3811; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3813 = 8'he5 == io_in_2 ? 8'h8c : _GEN_3812; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3814 = 8'he6 == io_in_2 ? 8'h97 : _GEN_3813; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3815 = 8'he7 == io_in_2 ? 8'h9e : _GEN_3814; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3816 = 8'he8 == io_in_2 ? 8'he9 : _GEN_3815; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3817 = 8'he9 == io_in_2 ? 8'he0 : _GEN_3816; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3818 = 8'hea == io_in_2 ? 8'hfb : _GEN_3817; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3819 = 8'heb == io_in_2 ? 8'hf2 : _GEN_3818; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3820 = 8'hec == io_in_2 ? 8'hcd : _GEN_3819; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3821 = 8'hed == io_in_2 ? 8'hc4 : _GEN_3820; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3822 = 8'hee == io_in_2 ? 8'hdf : _GEN_3821; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3823 = 8'hef == io_in_2 ? 8'hd6 : _GEN_3822; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3824 = 8'hf0 == io_in_2 ? 8'h31 : _GEN_3823; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3825 = 8'hf1 == io_in_2 ? 8'h38 : _GEN_3824; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3826 = 8'hf2 == io_in_2 ? 8'h23 : _GEN_3825; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3827 = 8'hf3 == io_in_2 ? 8'h2a : _GEN_3826; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3828 = 8'hf4 == io_in_2 ? 8'h15 : _GEN_3827; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3829 = 8'hf5 == io_in_2 ? 8'h1c : _GEN_3828; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3830 = 8'hf6 == io_in_2 ? 8'h7 : _GEN_3829; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3831 = 8'hf7 == io_in_2 ? 8'he : _GEN_3830; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3832 = 8'hf8 == io_in_2 ? 8'h79 : _GEN_3831; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3833 = 8'hf9 == io_in_2 ? 8'h70 : _GEN_3832; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3834 = 8'hfa == io_in_2 ? 8'h6b : _GEN_3833; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3835 = 8'hfb == io_in_2 ? 8'h62 : _GEN_3834; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3836 = 8'hfc == io_in_2 ? 8'h5d : _GEN_3835; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3837 = 8'hfd == io_in_2 ? 8'h54 : _GEN_3836; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3838 = 8'hfe == io_in_2 ? 8'h4f : _GEN_3837; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3839 = 8'hff == io_in_2 ? 8'h46 : _GEN_3838; // @[AES_PipelinedElasticBuffer.scala 594:50 AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _T_10 = _T_9 ^ _GEN_3839; // @[AES_PipelinedElasticBuffer.scala 594:50]
  wire [7:0] _GEN_3841 = 8'h1 == io_in_3 ? 8'he : 8'h0; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3842 = 8'h2 == io_in_3 ? 8'h1c : _GEN_3841; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3843 = 8'h3 == io_in_3 ? 8'h12 : _GEN_3842; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3844 = 8'h4 == io_in_3 ? 8'h38 : _GEN_3843; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3845 = 8'h5 == io_in_3 ? 8'h36 : _GEN_3844; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3846 = 8'h6 == io_in_3 ? 8'h24 : _GEN_3845; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3847 = 8'h7 == io_in_3 ? 8'h2a : _GEN_3846; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3848 = 8'h8 == io_in_3 ? 8'h70 : _GEN_3847; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3849 = 8'h9 == io_in_3 ? 8'h7e : _GEN_3848; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3850 = 8'ha == io_in_3 ? 8'h6c : _GEN_3849; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3851 = 8'hb == io_in_3 ? 8'h62 : _GEN_3850; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3852 = 8'hc == io_in_3 ? 8'h48 : _GEN_3851; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3853 = 8'hd == io_in_3 ? 8'h46 : _GEN_3852; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3854 = 8'he == io_in_3 ? 8'h54 : _GEN_3853; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3855 = 8'hf == io_in_3 ? 8'h5a : _GEN_3854; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3856 = 8'h10 == io_in_3 ? 8'he0 : _GEN_3855; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3857 = 8'h11 == io_in_3 ? 8'hee : _GEN_3856; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3858 = 8'h12 == io_in_3 ? 8'hfc : _GEN_3857; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3859 = 8'h13 == io_in_3 ? 8'hf2 : _GEN_3858; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3860 = 8'h14 == io_in_3 ? 8'hd8 : _GEN_3859; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3861 = 8'h15 == io_in_3 ? 8'hd6 : _GEN_3860; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3862 = 8'h16 == io_in_3 ? 8'hc4 : _GEN_3861; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3863 = 8'h17 == io_in_3 ? 8'hca : _GEN_3862; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3864 = 8'h18 == io_in_3 ? 8'h90 : _GEN_3863; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3865 = 8'h19 == io_in_3 ? 8'h9e : _GEN_3864; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3866 = 8'h1a == io_in_3 ? 8'h8c : _GEN_3865; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3867 = 8'h1b == io_in_3 ? 8'h82 : _GEN_3866; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3868 = 8'h1c == io_in_3 ? 8'ha8 : _GEN_3867; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3869 = 8'h1d == io_in_3 ? 8'ha6 : _GEN_3868; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3870 = 8'h1e == io_in_3 ? 8'hb4 : _GEN_3869; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3871 = 8'h1f == io_in_3 ? 8'hba : _GEN_3870; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3872 = 8'h20 == io_in_3 ? 8'hdb : _GEN_3871; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3873 = 8'h21 == io_in_3 ? 8'hd5 : _GEN_3872; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3874 = 8'h22 == io_in_3 ? 8'hc7 : _GEN_3873; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3875 = 8'h23 == io_in_3 ? 8'hc9 : _GEN_3874; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3876 = 8'h24 == io_in_3 ? 8'he3 : _GEN_3875; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3877 = 8'h25 == io_in_3 ? 8'hed : _GEN_3876; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3878 = 8'h26 == io_in_3 ? 8'hff : _GEN_3877; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3879 = 8'h27 == io_in_3 ? 8'hf1 : _GEN_3878; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3880 = 8'h28 == io_in_3 ? 8'hab : _GEN_3879; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3881 = 8'h29 == io_in_3 ? 8'ha5 : _GEN_3880; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3882 = 8'h2a == io_in_3 ? 8'hb7 : _GEN_3881; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3883 = 8'h2b == io_in_3 ? 8'hb9 : _GEN_3882; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3884 = 8'h2c == io_in_3 ? 8'h93 : _GEN_3883; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3885 = 8'h2d == io_in_3 ? 8'h9d : _GEN_3884; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3886 = 8'h2e == io_in_3 ? 8'h8f : _GEN_3885; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3887 = 8'h2f == io_in_3 ? 8'h81 : _GEN_3886; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3888 = 8'h30 == io_in_3 ? 8'h3b : _GEN_3887; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3889 = 8'h31 == io_in_3 ? 8'h35 : _GEN_3888; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3890 = 8'h32 == io_in_3 ? 8'h27 : _GEN_3889; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3891 = 8'h33 == io_in_3 ? 8'h29 : _GEN_3890; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3892 = 8'h34 == io_in_3 ? 8'h3 : _GEN_3891; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3893 = 8'h35 == io_in_3 ? 8'hd : _GEN_3892; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3894 = 8'h36 == io_in_3 ? 8'h1f : _GEN_3893; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3895 = 8'h37 == io_in_3 ? 8'h11 : _GEN_3894; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3896 = 8'h38 == io_in_3 ? 8'h4b : _GEN_3895; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3897 = 8'h39 == io_in_3 ? 8'h45 : _GEN_3896; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3898 = 8'h3a == io_in_3 ? 8'h57 : _GEN_3897; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3899 = 8'h3b == io_in_3 ? 8'h59 : _GEN_3898; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3900 = 8'h3c == io_in_3 ? 8'h73 : _GEN_3899; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3901 = 8'h3d == io_in_3 ? 8'h7d : _GEN_3900; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3902 = 8'h3e == io_in_3 ? 8'h6f : _GEN_3901; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3903 = 8'h3f == io_in_3 ? 8'h61 : _GEN_3902; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3904 = 8'h40 == io_in_3 ? 8'had : _GEN_3903; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3905 = 8'h41 == io_in_3 ? 8'ha3 : _GEN_3904; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3906 = 8'h42 == io_in_3 ? 8'hb1 : _GEN_3905; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3907 = 8'h43 == io_in_3 ? 8'hbf : _GEN_3906; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3908 = 8'h44 == io_in_3 ? 8'h95 : _GEN_3907; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3909 = 8'h45 == io_in_3 ? 8'h9b : _GEN_3908; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3910 = 8'h46 == io_in_3 ? 8'h89 : _GEN_3909; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3911 = 8'h47 == io_in_3 ? 8'h87 : _GEN_3910; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3912 = 8'h48 == io_in_3 ? 8'hdd : _GEN_3911; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3913 = 8'h49 == io_in_3 ? 8'hd3 : _GEN_3912; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3914 = 8'h4a == io_in_3 ? 8'hc1 : _GEN_3913; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3915 = 8'h4b == io_in_3 ? 8'hcf : _GEN_3914; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3916 = 8'h4c == io_in_3 ? 8'he5 : _GEN_3915; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3917 = 8'h4d == io_in_3 ? 8'heb : _GEN_3916; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3918 = 8'h4e == io_in_3 ? 8'hf9 : _GEN_3917; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3919 = 8'h4f == io_in_3 ? 8'hf7 : _GEN_3918; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3920 = 8'h50 == io_in_3 ? 8'h4d : _GEN_3919; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3921 = 8'h51 == io_in_3 ? 8'h43 : _GEN_3920; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3922 = 8'h52 == io_in_3 ? 8'h51 : _GEN_3921; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3923 = 8'h53 == io_in_3 ? 8'h5f : _GEN_3922; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3924 = 8'h54 == io_in_3 ? 8'h75 : _GEN_3923; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3925 = 8'h55 == io_in_3 ? 8'h7b : _GEN_3924; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3926 = 8'h56 == io_in_3 ? 8'h69 : _GEN_3925; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3927 = 8'h57 == io_in_3 ? 8'h67 : _GEN_3926; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3928 = 8'h58 == io_in_3 ? 8'h3d : _GEN_3927; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3929 = 8'h59 == io_in_3 ? 8'h33 : _GEN_3928; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3930 = 8'h5a == io_in_3 ? 8'h21 : _GEN_3929; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3931 = 8'h5b == io_in_3 ? 8'h2f : _GEN_3930; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3932 = 8'h5c == io_in_3 ? 8'h5 : _GEN_3931; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3933 = 8'h5d == io_in_3 ? 8'hb : _GEN_3932; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3934 = 8'h5e == io_in_3 ? 8'h19 : _GEN_3933; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3935 = 8'h5f == io_in_3 ? 8'h17 : _GEN_3934; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3936 = 8'h60 == io_in_3 ? 8'h76 : _GEN_3935; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3937 = 8'h61 == io_in_3 ? 8'h78 : _GEN_3936; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3938 = 8'h62 == io_in_3 ? 8'h6a : _GEN_3937; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3939 = 8'h63 == io_in_3 ? 8'h64 : _GEN_3938; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3940 = 8'h64 == io_in_3 ? 8'h4e : _GEN_3939; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3941 = 8'h65 == io_in_3 ? 8'h40 : _GEN_3940; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3942 = 8'h66 == io_in_3 ? 8'h52 : _GEN_3941; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3943 = 8'h67 == io_in_3 ? 8'h5c : _GEN_3942; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3944 = 8'h68 == io_in_3 ? 8'h6 : _GEN_3943; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3945 = 8'h69 == io_in_3 ? 8'h8 : _GEN_3944; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3946 = 8'h6a == io_in_3 ? 8'h1a : _GEN_3945; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3947 = 8'h6b == io_in_3 ? 8'h14 : _GEN_3946; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3948 = 8'h6c == io_in_3 ? 8'h3e : _GEN_3947; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3949 = 8'h6d == io_in_3 ? 8'h30 : _GEN_3948; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3950 = 8'h6e == io_in_3 ? 8'h22 : _GEN_3949; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3951 = 8'h6f == io_in_3 ? 8'h2c : _GEN_3950; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3952 = 8'h70 == io_in_3 ? 8'h96 : _GEN_3951; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3953 = 8'h71 == io_in_3 ? 8'h98 : _GEN_3952; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3954 = 8'h72 == io_in_3 ? 8'h8a : _GEN_3953; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3955 = 8'h73 == io_in_3 ? 8'h84 : _GEN_3954; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3956 = 8'h74 == io_in_3 ? 8'hae : _GEN_3955; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3957 = 8'h75 == io_in_3 ? 8'ha0 : _GEN_3956; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3958 = 8'h76 == io_in_3 ? 8'hb2 : _GEN_3957; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3959 = 8'h77 == io_in_3 ? 8'hbc : _GEN_3958; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3960 = 8'h78 == io_in_3 ? 8'he6 : _GEN_3959; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3961 = 8'h79 == io_in_3 ? 8'he8 : _GEN_3960; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3962 = 8'h7a == io_in_3 ? 8'hfa : _GEN_3961; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3963 = 8'h7b == io_in_3 ? 8'hf4 : _GEN_3962; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3964 = 8'h7c == io_in_3 ? 8'hde : _GEN_3963; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3965 = 8'h7d == io_in_3 ? 8'hd0 : _GEN_3964; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3966 = 8'h7e == io_in_3 ? 8'hc2 : _GEN_3965; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3967 = 8'h7f == io_in_3 ? 8'hcc : _GEN_3966; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3968 = 8'h80 == io_in_3 ? 8'h41 : _GEN_3967; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3969 = 8'h81 == io_in_3 ? 8'h4f : _GEN_3968; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3970 = 8'h82 == io_in_3 ? 8'h5d : _GEN_3969; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3971 = 8'h83 == io_in_3 ? 8'h53 : _GEN_3970; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3972 = 8'h84 == io_in_3 ? 8'h79 : _GEN_3971; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3973 = 8'h85 == io_in_3 ? 8'h77 : _GEN_3972; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3974 = 8'h86 == io_in_3 ? 8'h65 : _GEN_3973; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3975 = 8'h87 == io_in_3 ? 8'h6b : _GEN_3974; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3976 = 8'h88 == io_in_3 ? 8'h31 : _GEN_3975; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3977 = 8'h89 == io_in_3 ? 8'h3f : _GEN_3976; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3978 = 8'h8a == io_in_3 ? 8'h2d : _GEN_3977; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3979 = 8'h8b == io_in_3 ? 8'h23 : _GEN_3978; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3980 = 8'h8c == io_in_3 ? 8'h9 : _GEN_3979; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3981 = 8'h8d == io_in_3 ? 8'h7 : _GEN_3980; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3982 = 8'h8e == io_in_3 ? 8'h15 : _GEN_3981; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3983 = 8'h8f == io_in_3 ? 8'h1b : _GEN_3982; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3984 = 8'h90 == io_in_3 ? 8'ha1 : _GEN_3983; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3985 = 8'h91 == io_in_3 ? 8'haf : _GEN_3984; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3986 = 8'h92 == io_in_3 ? 8'hbd : _GEN_3985; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3987 = 8'h93 == io_in_3 ? 8'hb3 : _GEN_3986; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3988 = 8'h94 == io_in_3 ? 8'h99 : _GEN_3987; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3989 = 8'h95 == io_in_3 ? 8'h97 : _GEN_3988; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3990 = 8'h96 == io_in_3 ? 8'h85 : _GEN_3989; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3991 = 8'h97 == io_in_3 ? 8'h8b : _GEN_3990; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3992 = 8'h98 == io_in_3 ? 8'hd1 : _GEN_3991; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3993 = 8'h99 == io_in_3 ? 8'hdf : _GEN_3992; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3994 = 8'h9a == io_in_3 ? 8'hcd : _GEN_3993; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3995 = 8'h9b == io_in_3 ? 8'hc3 : _GEN_3994; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3996 = 8'h9c == io_in_3 ? 8'he9 : _GEN_3995; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3997 = 8'h9d == io_in_3 ? 8'he7 : _GEN_3996; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3998 = 8'h9e == io_in_3 ? 8'hf5 : _GEN_3997; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_3999 = 8'h9f == io_in_3 ? 8'hfb : _GEN_3998; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4000 = 8'ha0 == io_in_3 ? 8'h9a : _GEN_3999; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4001 = 8'ha1 == io_in_3 ? 8'h94 : _GEN_4000; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4002 = 8'ha2 == io_in_3 ? 8'h86 : _GEN_4001; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4003 = 8'ha3 == io_in_3 ? 8'h88 : _GEN_4002; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4004 = 8'ha4 == io_in_3 ? 8'ha2 : _GEN_4003; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4005 = 8'ha5 == io_in_3 ? 8'hac : _GEN_4004; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4006 = 8'ha6 == io_in_3 ? 8'hbe : _GEN_4005; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4007 = 8'ha7 == io_in_3 ? 8'hb0 : _GEN_4006; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4008 = 8'ha8 == io_in_3 ? 8'hea : _GEN_4007; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4009 = 8'ha9 == io_in_3 ? 8'he4 : _GEN_4008; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4010 = 8'haa == io_in_3 ? 8'hf6 : _GEN_4009; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4011 = 8'hab == io_in_3 ? 8'hf8 : _GEN_4010; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4012 = 8'hac == io_in_3 ? 8'hd2 : _GEN_4011; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4013 = 8'had == io_in_3 ? 8'hdc : _GEN_4012; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4014 = 8'hae == io_in_3 ? 8'hce : _GEN_4013; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4015 = 8'haf == io_in_3 ? 8'hc0 : _GEN_4014; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4016 = 8'hb0 == io_in_3 ? 8'h7a : _GEN_4015; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4017 = 8'hb1 == io_in_3 ? 8'h74 : _GEN_4016; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4018 = 8'hb2 == io_in_3 ? 8'h66 : _GEN_4017; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4019 = 8'hb3 == io_in_3 ? 8'h68 : _GEN_4018; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4020 = 8'hb4 == io_in_3 ? 8'h42 : _GEN_4019; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4021 = 8'hb5 == io_in_3 ? 8'h4c : _GEN_4020; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4022 = 8'hb6 == io_in_3 ? 8'h5e : _GEN_4021; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4023 = 8'hb7 == io_in_3 ? 8'h50 : _GEN_4022; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4024 = 8'hb8 == io_in_3 ? 8'ha : _GEN_4023; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4025 = 8'hb9 == io_in_3 ? 8'h4 : _GEN_4024; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4026 = 8'hba == io_in_3 ? 8'h16 : _GEN_4025; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4027 = 8'hbb == io_in_3 ? 8'h18 : _GEN_4026; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4028 = 8'hbc == io_in_3 ? 8'h32 : _GEN_4027; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4029 = 8'hbd == io_in_3 ? 8'h3c : _GEN_4028; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4030 = 8'hbe == io_in_3 ? 8'h2e : _GEN_4029; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4031 = 8'hbf == io_in_3 ? 8'h20 : _GEN_4030; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4032 = 8'hc0 == io_in_3 ? 8'hec : _GEN_4031; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4033 = 8'hc1 == io_in_3 ? 8'he2 : _GEN_4032; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4034 = 8'hc2 == io_in_3 ? 8'hf0 : _GEN_4033; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4035 = 8'hc3 == io_in_3 ? 8'hfe : _GEN_4034; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4036 = 8'hc4 == io_in_3 ? 8'hd4 : _GEN_4035; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4037 = 8'hc5 == io_in_3 ? 8'hda : _GEN_4036; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4038 = 8'hc6 == io_in_3 ? 8'hc8 : _GEN_4037; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4039 = 8'hc7 == io_in_3 ? 8'hc6 : _GEN_4038; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4040 = 8'hc8 == io_in_3 ? 8'h9c : _GEN_4039; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4041 = 8'hc9 == io_in_3 ? 8'h92 : _GEN_4040; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4042 = 8'hca == io_in_3 ? 8'h80 : _GEN_4041; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4043 = 8'hcb == io_in_3 ? 8'h8e : _GEN_4042; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4044 = 8'hcc == io_in_3 ? 8'ha4 : _GEN_4043; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4045 = 8'hcd == io_in_3 ? 8'haa : _GEN_4044; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4046 = 8'hce == io_in_3 ? 8'hb8 : _GEN_4045; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4047 = 8'hcf == io_in_3 ? 8'hb6 : _GEN_4046; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4048 = 8'hd0 == io_in_3 ? 8'hc : _GEN_4047; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4049 = 8'hd1 == io_in_3 ? 8'h2 : _GEN_4048; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4050 = 8'hd2 == io_in_3 ? 8'h10 : _GEN_4049; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4051 = 8'hd3 == io_in_3 ? 8'h1e : _GEN_4050; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4052 = 8'hd4 == io_in_3 ? 8'h34 : _GEN_4051; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4053 = 8'hd5 == io_in_3 ? 8'h3a : _GEN_4052; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4054 = 8'hd6 == io_in_3 ? 8'h28 : _GEN_4053; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4055 = 8'hd7 == io_in_3 ? 8'h26 : _GEN_4054; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4056 = 8'hd8 == io_in_3 ? 8'h7c : _GEN_4055; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4057 = 8'hd9 == io_in_3 ? 8'h72 : _GEN_4056; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4058 = 8'hda == io_in_3 ? 8'h60 : _GEN_4057; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4059 = 8'hdb == io_in_3 ? 8'h6e : _GEN_4058; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4060 = 8'hdc == io_in_3 ? 8'h44 : _GEN_4059; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4061 = 8'hdd == io_in_3 ? 8'h4a : _GEN_4060; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4062 = 8'hde == io_in_3 ? 8'h58 : _GEN_4061; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4063 = 8'hdf == io_in_3 ? 8'h56 : _GEN_4062; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4064 = 8'he0 == io_in_3 ? 8'h37 : _GEN_4063; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4065 = 8'he1 == io_in_3 ? 8'h39 : _GEN_4064; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4066 = 8'he2 == io_in_3 ? 8'h2b : _GEN_4065; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4067 = 8'he3 == io_in_3 ? 8'h25 : _GEN_4066; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4068 = 8'he4 == io_in_3 ? 8'hf : _GEN_4067; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4069 = 8'he5 == io_in_3 ? 8'h1 : _GEN_4068; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4070 = 8'he6 == io_in_3 ? 8'h13 : _GEN_4069; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4071 = 8'he7 == io_in_3 ? 8'h1d : _GEN_4070; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4072 = 8'he8 == io_in_3 ? 8'h47 : _GEN_4071; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4073 = 8'he9 == io_in_3 ? 8'h49 : _GEN_4072; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4074 = 8'hea == io_in_3 ? 8'h5b : _GEN_4073; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4075 = 8'heb == io_in_3 ? 8'h55 : _GEN_4074; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4076 = 8'hec == io_in_3 ? 8'h7f : _GEN_4075; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4077 = 8'hed == io_in_3 ? 8'h71 : _GEN_4076; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4078 = 8'hee == io_in_3 ? 8'h63 : _GEN_4077; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4079 = 8'hef == io_in_3 ? 8'h6d : _GEN_4078; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4080 = 8'hf0 == io_in_3 ? 8'hd7 : _GEN_4079; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4081 = 8'hf1 == io_in_3 ? 8'hd9 : _GEN_4080; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4082 = 8'hf2 == io_in_3 ? 8'hcb : _GEN_4081; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4083 = 8'hf3 == io_in_3 ? 8'hc5 : _GEN_4082; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4084 = 8'hf4 == io_in_3 ? 8'hef : _GEN_4083; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4085 = 8'hf5 == io_in_3 ? 8'he1 : _GEN_4084; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4086 = 8'hf6 == io_in_3 ? 8'hf3 : _GEN_4085; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4087 = 8'hf7 == io_in_3 ? 8'hfd : _GEN_4086; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4088 = 8'hf8 == io_in_3 ? 8'ha7 : _GEN_4087; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4089 = 8'hf9 == io_in_3 ? 8'ha9 : _GEN_4088; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4090 = 8'hfa == io_in_3 ? 8'hbb : _GEN_4089; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4091 = 8'hfb == io_in_3 ? 8'hb5 : _GEN_4090; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4092 = 8'hfc == io_in_3 ? 8'h9f : _GEN_4091; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4093 = 8'hfd == io_in_3 ? 8'h91 : _GEN_4092; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4094 = 8'hfe == io_in_3 ? 8'h83 : _GEN_4093; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  wire [7:0] _GEN_4095 = 8'hff == io_in_3 ? 8'h8d : _GEN_4094; // @[AES_PipelinedElasticBuffer.scala 594:67 AES_PipelinedElasticBuffer.scala 594:67]
  assign io_out_0 = _T_1 ^ _GEN_1023; // @[AES_PipelinedElasticBuffer.scala 591:68]
  assign io_out_1 = _T_4 ^ _GEN_2047; // @[AES_PipelinedElasticBuffer.scala 592:67]
  assign io_out_2 = _T_7 ^ _GEN_3071; // @[AES_PipelinedElasticBuffer.scala 593:67]
  assign io_out_3 = _T_10 ^ _GEN_4095; // @[AES_PipelinedElasticBuffer.scala 594:67]
endmodule
module AES_InvMixColumns(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3
);
  wire [7:0] PEs_0_io_in_0; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_0_io_in_1; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_0_io_in_2; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_0_io_in_3; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_0_io_out_0; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_0_io_out_1; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_0_io_out_2; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_0_io_out_3; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_1_io_in_0; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_1_io_in_1; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_1_io_in_2; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_1_io_in_3; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_1_io_out_0; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_1_io_out_1; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_1_io_out_2; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_1_io_out_3; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_2_io_in_0; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_2_io_in_1; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_2_io_in_2; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_2_io_in_3; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_2_io_out_0; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_2_io_out_1; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_2_io_out_2; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_2_io_out_3; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_3_io_in_0; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_3_io_in_1; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_3_io_in_2; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_3_io_in_3; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_3_io_out_0; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_3_io_out_1; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_3_io_out_2; // @[AES_PipelinedElasticBuffer.scala 397:20]
  wire [7:0] PEs_3_io_out_3; // @[AES_PipelinedElasticBuffer.scala 397:20]
  AES_InvMixColumn PEs_0 ( // @[AES_PipelinedElasticBuffer.scala 397:20]
    .io_in_0(PEs_0_io_in_0),
    .io_in_1(PEs_0_io_in_1),
    .io_in_2(PEs_0_io_in_2),
    .io_in_3(PEs_0_io_in_3),
    .io_out_0(PEs_0_io_out_0),
    .io_out_1(PEs_0_io_out_1),
    .io_out_2(PEs_0_io_out_2),
    .io_out_3(PEs_0_io_out_3)
  );
  AES_InvMixColumn PEs_1 ( // @[AES_PipelinedElasticBuffer.scala 397:20]
    .io_in_0(PEs_1_io_in_0),
    .io_in_1(PEs_1_io_in_1),
    .io_in_2(PEs_1_io_in_2),
    .io_in_3(PEs_1_io_in_3),
    .io_out_0(PEs_1_io_out_0),
    .io_out_1(PEs_1_io_out_1),
    .io_out_2(PEs_1_io_out_2),
    .io_out_3(PEs_1_io_out_3)
  );
  AES_InvMixColumn PEs_2 ( // @[AES_PipelinedElasticBuffer.scala 397:20]
    .io_in_0(PEs_2_io_in_0),
    .io_in_1(PEs_2_io_in_1),
    .io_in_2(PEs_2_io_in_2),
    .io_in_3(PEs_2_io_in_3),
    .io_out_0(PEs_2_io_out_0),
    .io_out_1(PEs_2_io_out_1),
    .io_out_2(PEs_2_io_out_2),
    .io_out_3(PEs_2_io_out_3)
  );
  AES_InvMixColumn PEs_3 ( // @[AES_PipelinedElasticBuffer.scala 397:20]
    .io_in_0(PEs_3_io_in_0),
    .io_in_1(PEs_3_io_in_1),
    .io_in_2(PEs_3_io_in_2),
    .io_in_3(PEs_3_io_in_3),
    .io_out_0(PEs_3_io_out_0),
    .io_out_1(PEs_3_io_out_1),
    .io_out_2(PEs_3_io_out_2),
    .io_out_3(PEs_3_io_out_3)
  );
  assign io_out_state_0_0 = PEs_0_io_out_0; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_0_1 = PEs_0_io_out_1; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_0_2 = PEs_0_io_out_2; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_0_3 = PEs_0_io_out_3; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_1_0 = PEs_1_io_out_0; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_1_1 = PEs_1_io_out_1; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_1_2 = PEs_1_io_out_2; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_1_3 = PEs_1_io_out_3; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_2_0 = PEs_2_io_out_0; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_2_1 = PEs_2_io_out_1; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_2_2 = PEs_2_io_out_2; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_2_3 = PEs_2_io_out_3; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_3_0 = PEs_3_io_out_0; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_3_1 = PEs_3_io_out_1; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_3_2 = PEs_3_io_out_2; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign io_out_state_3_3 = PEs_3_io_out_3; // @[AES_PipelinedElasticBuffer.scala 404:21]
  assign PEs_0_io_in_0 = io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_0_io_in_1 = io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_0_io_in_2 = io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_0_io_in_3 = io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_1_io_in_0 = io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_1_io_in_1 = io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_1_io_in_2 = io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_1_io_in_3 = io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_2_io_in_0 = io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_2_io_in_1 = io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_2_io_in_2 = io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_2_io_in_3 = io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_3_io_in_0 = io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_3_io_in_1 = io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_3_io_in_2 = io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 403:18]
  assign PEs_3_io_in_3 = io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 403:18]
endmodule
module AES_InvShiftRows(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3
);
  assign io_out_state_0_0 = io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 634:22]
  assign io_out_state_0_1 = io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 639:22]
  assign io_out_state_0_2 = io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 644:22]
  assign io_out_state_0_3 = io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 649:22]
  assign io_out_state_1_0 = io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 635:22]
  assign io_out_state_1_1 = io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 640:22]
  assign io_out_state_1_2 = io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 645:22]
  assign io_out_state_1_3 = io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 650:22]
  assign io_out_state_2_0 = io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 636:22]
  assign io_out_state_2_1 = io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 641:22]
  assign io_out_state_2_2 = io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 646:22]
  assign io_out_state_2_3 = io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 651:22]
  assign io_out_state_3_0 = io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 637:22]
  assign io_out_state_3_1 = io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 642:22]
  assign io_out_state_3_2 = io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 647:22]
  assign io_out_state_3_3 = io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 652:22]
endmodule
module AES_InvS(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _GEN_1 = 4'h0 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h9 : 8'h52; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_2 = 4'h0 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h6a : _GEN_1; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_3 = 4'h0 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hd5 : _GEN_2; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_4 = 4'h0 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h30 : _GEN_3; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_5 = 4'h0 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h36 : _GEN_4; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_6 = 4'h0 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'ha5 : _GEN_5; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_7 = 4'h0 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h38 : _GEN_6; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_8 = 4'h0 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hbf : _GEN_7; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_9 = 4'h0 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h40 : _GEN_8; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_10 = 4'h0 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'ha3 : _GEN_9; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_11 = 4'h0 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h9e : _GEN_10; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_12 = 4'h0 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h81 : _GEN_11; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_13 = 4'h0 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hf3 : _GEN_12; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_14 = 4'h0 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hd7 : _GEN_13; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_15 = 4'h0 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hfb : _GEN_14; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_16 = 4'h1 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h7c : _GEN_15; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_17 = 4'h1 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'he3 : _GEN_16; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_18 = 4'h1 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h39 : _GEN_17; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_19 = 4'h1 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h82 : _GEN_18; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_20 = 4'h1 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h9b : _GEN_19; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_21 = 4'h1 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h2f : _GEN_20; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_22 = 4'h1 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hff : _GEN_21; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_23 = 4'h1 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h87 : _GEN_22; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_24 = 4'h1 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h34 : _GEN_23; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_25 = 4'h1 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h8e : _GEN_24; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_26 = 4'h1 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h43 : _GEN_25; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_27 = 4'h1 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h44 : _GEN_26; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_28 = 4'h1 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hc4 : _GEN_27; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_29 = 4'h1 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hde : _GEN_28; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_30 = 4'h1 == io_in[7:4] & 4'he == io_in[3:0] ? 8'he9 : _GEN_29; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_31 = 4'h1 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hcb : _GEN_30; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_32 = 4'h2 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h54 : _GEN_31; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_33 = 4'h2 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h7b : _GEN_32; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_34 = 4'h2 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h94 : _GEN_33; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_35 = 4'h2 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h32 : _GEN_34; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_36 = 4'h2 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'ha6 : _GEN_35; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_37 = 4'h2 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hc2 : _GEN_36; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_38 = 4'h2 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h23 : _GEN_37; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_39 = 4'h2 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h3d : _GEN_38; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_40 = 4'h2 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hee : _GEN_39; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_41 = 4'h2 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h4c : _GEN_40; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_42 = 4'h2 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h95 : _GEN_41; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_43 = 4'h2 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hb : _GEN_42; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_44 = 4'h2 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h42 : _GEN_43; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_45 = 4'h2 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hfa : _GEN_44; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_46 = 4'h2 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hc3 : _GEN_45; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_47 = 4'h2 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h4e : _GEN_46; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_48 = 4'h3 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h8 : _GEN_47; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_49 = 4'h3 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h2e : _GEN_48; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_50 = 4'h3 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'ha1 : _GEN_49; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_51 = 4'h3 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h66 : _GEN_50; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_52 = 4'h3 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h28 : _GEN_51; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_53 = 4'h3 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hd9 : _GEN_52; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_54 = 4'h3 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h24 : _GEN_53; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_55 = 4'h3 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hb2 : _GEN_54; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_56 = 4'h3 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h76 : _GEN_55; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_57 = 4'h3 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h5b : _GEN_56; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_58 = 4'h3 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'ha2 : _GEN_57; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_59 = 4'h3 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h49 : _GEN_58; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_60 = 4'h3 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h6d : _GEN_59; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_61 = 4'h3 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h8b : _GEN_60; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_62 = 4'h3 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hd1 : _GEN_61; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_63 = 4'h3 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h25 : _GEN_62; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_64 = 4'h4 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h72 : _GEN_63; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_65 = 4'h4 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hf8 : _GEN_64; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_66 = 4'h4 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'hf6 : _GEN_65; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_67 = 4'h4 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h64 : _GEN_66; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_68 = 4'h4 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h86 : _GEN_67; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_69 = 4'h4 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h68 : _GEN_68; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_70 = 4'h4 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h98 : _GEN_69; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_71 = 4'h4 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h16 : _GEN_70; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_72 = 4'h4 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hd4 : _GEN_71; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_73 = 4'h4 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'ha4 : _GEN_72; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_74 = 4'h4 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h5c : _GEN_73; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_75 = 4'h4 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hcc : _GEN_74; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_76 = 4'h4 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h5d : _GEN_75; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_77 = 4'h4 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h65 : _GEN_76; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_78 = 4'h4 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hb6 : _GEN_77; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_79 = 4'h4 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h92 : _GEN_78; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_80 = 4'h5 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h6c : _GEN_79; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_81 = 4'h5 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h70 : _GEN_80; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_82 = 4'h5 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h48 : _GEN_81; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_83 = 4'h5 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h50 : _GEN_82; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_84 = 4'h5 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hfd : _GEN_83; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_85 = 4'h5 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hed : _GEN_84; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_86 = 4'h5 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hb9 : _GEN_85; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_87 = 4'h5 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hda : _GEN_86; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_88 = 4'h5 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h5e : _GEN_87; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_89 = 4'h5 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h15 : _GEN_88; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_90 = 4'h5 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h46 : _GEN_89; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_91 = 4'h5 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h57 : _GEN_90; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_92 = 4'h5 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'ha7 : _GEN_91; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_93 = 4'h5 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h8d : _GEN_92; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_94 = 4'h5 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h9d : _GEN_93; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_95 = 4'h5 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h84 : _GEN_94; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_96 = 4'h6 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h90 : _GEN_95; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_97 = 4'h6 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hd8 : _GEN_96; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_98 = 4'h6 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'hab : _GEN_97; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_99 = 4'h6 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h0 : _GEN_98; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_100 = 4'h6 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h8c : _GEN_99; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_101 = 4'h6 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hbc : _GEN_100; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_102 = 4'h6 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hd3 : _GEN_101; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_103 = 4'h6 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'ha : _GEN_102; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_104 = 4'h6 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hf7 : _GEN_103; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_105 = 4'h6 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'he4 : _GEN_104; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_106 = 4'h6 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h58 : _GEN_105; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_107 = 4'h6 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h5 : _GEN_106; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_108 = 4'h6 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hb8 : _GEN_107; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_109 = 4'h6 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hb3 : _GEN_108; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_110 = 4'h6 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h45 : _GEN_109; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_111 = 4'h6 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h6 : _GEN_110; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_112 = 4'h7 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hd0 : _GEN_111; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_113 = 4'h7 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h2c : _GEN_112; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_114 = 4'h7 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h1e : _GEN_113; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_115 = 4'h7 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h8f : _GEN_114; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_116 = 4'h7 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hca : _GEN_115; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_117 = 4'h7 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h3f : _GEN_116; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_118 = 4'h7 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hf : _GEN_117; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_119 = 4'h7 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h2 : _GEN_118; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_120 = 4'h7 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hc1 : _GEN_119; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_121 = 4'h7 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'haf : _GEN_120; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_122 = 4'h7 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hbd : _GEN_121; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_123 = 4'h7 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h3 : _GEN_122; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_124 = 4'h7 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h1 : _GEN_123; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_125 = 4'h7 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h13 : _GEN_124; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_126 = 4'h7 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h8a : _GEN_125; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_127 = 4'h7 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h6b : _GEN_126; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_128 = 4'h8 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h3a : _GEN_127; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_129 = 4'h8 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h91 : _GEN_128; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_130 = 4'h8 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h11 : _GEN_129; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_131 = 4'h8 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h41 : _GEN_130; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_132 = 4'h8 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h4f : _GEN_131; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_133 = 4'h8 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h67 : _GEN_132; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_134 = 4'h8 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hdc : _GEN_133; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_135 = 4'h8 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hea : _GEN_134; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_136 = 4'h8 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h97 : _GEN_135; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_137 = 4'h8 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hf2 : _GEN_136; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_138 = 4'h8 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hcf : _GEN_137; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_139 = 4'h8 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hce : _GEN_138; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_140 = 4'h8 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hf0 : _GEN_139; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_141 = 4'h8 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hb4 : _GEN_140; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_142 = 4'h8 == io_in[7:4] & 4'he == io_in[3:0] ? 8'he6 : _GEN_141; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_143 = 4'h8 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h73 : _GEN_142; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_144 = 4'h9 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h96 : _GEN_143; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_145 = 4'h9 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hac : _GEN_144; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_146 = 4'h9 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h74 : _GEN_145; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_147 = 4'h9 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h22 : _GEN_146; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_148 = 4'h9 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'he7 : _GEN_147; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_149 = 4'h9 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'had : _GEN_148; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_150 = 4'h9 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h35 : _GEN_149; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_151 = 4'h9 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h85 : _GEN_150; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_152 = 4'h9 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'he2 : _GEN_151; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_153 = 4'h9 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hf9 : _GEN_152; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_154 = 4'h9 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h37 : _GEN_153; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_155 = 4'h9 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'he8 : _GEN_154; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_156 = 4'h9 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h1c : _GEN_155; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_157 = 4'h9 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h75 : _GEN_156; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_158 = 4'h9 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hdf : _GEN_157; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_159 = 4'h9 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h6e : _GEN_158; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_160 = 4'ha == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h47 : _GEN_159; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_161 = 4'ha == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hf1 : _GEN_160; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_162 = 4'ha == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h1a : _GEN_161; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_163 = 4'ha == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h71 : _GEN_162; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_164 = 4'ha == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h1d : _GEN_163; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_165 = 4'ha == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h29 : _GEN_164; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_166 = 4'ha == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hc5 : _GEN_165; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_167 = 4'ha == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h89 : _GEN_166; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_168 = 4'ha == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h6f : _GEN_167; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_169 = 4'ha == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hb7 : _GEN_168; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_170 = 4'ha == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h62 : _GEN_169; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_171 = 4'ha == io_in[7:4] & 4'hb == io_in[3:0] ? 8'he : _GEN_170; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_172 = 4'ha == io_in[7:4] & 4'hc == io_in[3:0] ? 8'haa : _GEN_171; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_173 = 4'ha == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h18 : _GEN_172; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_174 = 4'ha == io_in[7:4] & 4'he == io_in[3:0] ? 8'hbe : _GEN_173; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_175 = 4'ha == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h1b : _GEN_174; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_176 = 4'hb == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hfc : _GEN_175; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_177 = 4'hb == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h56 : _GEN_176; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_178 = 4'hb == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h3e : _GEN_177; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_179 = 4'hb == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h4b : _GEN_178; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_180 = 4'hb == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hc6 : _GEN_179; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_181 = 4'hb == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hd2 : _GEN_180; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_182 = 4'hb == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h79 : _GEN_181; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_183 = 4'hb == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h20 : _GEN_182; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_184 = 4'hb == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h9a : _GEN_183; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_185 = 4'hb == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hdb : _GEN_184; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_186 = 4'hb == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hc0 : _GEN_185; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_187 = 4'hb == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hfe : _GEN_186; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_188 = 4'hb == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h78 : _GEN_187; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_189 = 4'hb == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hcd : _GEN_188; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_190 = 4'hb == io_in[7:4] & 4'he == io_in[3:0] ? 8'h5a : _GEN_189; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_191 = 4'hb == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hf4 : _GEN_190; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_192 = 4'hc == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h1f : _GEN_191; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_193 = 4'hc == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hdd : _GEN_192; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_194 = 4'hc == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'ha8 : _GEN_193; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_195 = 4'hc == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h33 : _GEN_194; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_196 = 4'hc == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h88 : _GEN_195; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_197 = 4'hc == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h7 : _GEN_196; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_198 = 4'hc == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hc7 : _GEN_197; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_199 = 4'hc == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h31 : _GEN_198; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_200 = 4'hc == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hb1 : _GEN_199; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_201 = 4'hc == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h12 : _GEN_200; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_202 = 4'hc == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h10 : _GEN_201; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_203 = 4'hc == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h59 : _GEN_202; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_204 = 4'hc == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h27 : _GEN_203; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_205 = 4'hc == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h80 : _GEN_204; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_206 = 4'hc == io_in[7:4] & 4'he == io_in[3:0] ? 8'hec : _GEN_205; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_207 = 4'hc == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h5f : _GEN_206; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_208 = 4'hd == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h60 : _GEN_207; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_209 = 4'hd == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h51 : _GEN_208; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_210 = 4'hd == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h7f : _GEN_209; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_211 = 4'hd == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'ha9 : _GEN_210; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_212 = 4'hd == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h19 : _GEN_211; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_213 = 4'hd == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hb5 : _GEN_212; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_214 = 4'hd == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h4a : _GEN_213; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_215 = 4'hd == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hd : _GEN_214; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_216 = 4'hd == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h2d : _GEN_215; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_217 = 4'hd == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'he5 : _GEN_216; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_218 = 4'hd == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h7a : _GEN_217; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_219 = 4'hd == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h9f : _GEN_218; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_220 = 4'hd == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h93 : _GEN_219; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_221 = 4'hd == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hc9 : _GEN_220; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_222 = 4'hd == io_in[7:4] & 4'he == io_in[3:0] ? 8'h9c : _GEN_221; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_223 = 4'hd == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hef : _GEN_222; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_224 = 4'he == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'ha0 : _GEN_223; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_225 = 4'he == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'he0 : _GEN_224; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_226 = 4'he == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h3b : _GEN_225; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_227 = 4'he == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h4d : _GEN_226; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_228 = 4'he == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hae : _GEN_227; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_229 = 4'he == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h2a : _GEN_228; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_230 = 4'he == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hf5 : _GEN_229; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_231 = 4'he == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hb0 : _GEN_230; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_232 = 4'he == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hc8 : _GEN_231; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_233 = 4'he == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'heb : _GEN_232; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_234 = 4'he == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hbb : _GEN_233; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_235 = 4'he == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h3c : _GEN_234; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_236 = 4'he == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h83 : _GEN_235; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_237 = 4'he == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h53 : _GEN_236; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_238 = 4'he == io_in[7:4] & 4'he == io_in[3:0] ? 8'h99 : _GEN_237; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_239 = 4'he == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h61 : _GEN_238; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_240 = 4'hf == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h17 : _GEN_239; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_241 = 4'hf == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h2b : _GEN_240; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_242 = 4'hf == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h4 : _GEN_241; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_243 = 4'hf == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h7e : _GEN_242; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_244 = 4'hf == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hba : _GEN_243; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_245 = 4'hf == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h77 : _GEN_244; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_246 = 4'hf == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hd6 : _GEN_245; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_247 = 4'hf == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h26 : _GEN_246; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_248 = 4'hf == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'he1 : _GEN_247; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_249 = 4'hf == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h69 : _GEN_248; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_250 = 4'hf == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h14 : _GEN_249; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_251 = 4'hf == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h63 : _GEN_250; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_252 = 4'hf == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h55 : _GEN_251; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_253 = 4'hf == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h21 : _GEN_252; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  wire [7:0] _GEN_254 = 4'hf == io_in[7:4] & 4'he == io_in[3:0] ? 8'hc : _GEN_253; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
  assign io_out = 4'hf == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h7d : _GEN_254; // @[AES_PipelinedElasticBuffer.scala 784:10 AES_PipelinedElasticBuffer.scala 784:10]
endmodule
module AES_InvSubBytes(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3
);
  wire [7:0] invPEs_0_0_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_0_0_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_0_1_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_0_1_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_0_2_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_0_2_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_0_3_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_0_3_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_1_0_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_1_0_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_1_1_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_1_1_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_1_2_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_1_2_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_1_3_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_1_3_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_2_0_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_2_0_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_2_1_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_2_1_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_2_2_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_2_2_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_2_3_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_2_3_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_3_0_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_3_0_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_3_1_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_3_1_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_3_2_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_3_2_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_3_3_io_in; // @[AES_PipelinedElasticBuffer.scala 689:22]
  wire [7:0] invPEs_3_3_io_out; // @[AES_PipelinedElasticBuffer.scala 689:22]
  AES_InvS invPEs_0_0 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_0_0_io_in),
    .io_out(invPEs_0_0_io_out)
  );
  AES_InvS invPEs_0_1 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_0_1_io_in),
    .io_out(invPEs_0_1_io_out)
  );
  AES_InvS invPEs_0_2 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_0_2_io_in),
    .io_out(invPEs_0_2_io_out)
  );
  AES_InvS invPEs_0_3 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_0_3_io_in),
    .io_out(invPEs_0_3_io_out)
  );
  AES_InvS invPEs_1_0 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_1_0_io_in),
    .io_out(invPEs_1_0_io_out)
  );
  AES_InvS invPEs_1_1 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_1_1_io_in),
    .io_out(invPEs_1_1_io_out)
  );
  AES_InvS invPEs_1_2 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_1_2_io_in),
    .io_out(invPEs_1_2_io_out)
  );
  AES_InvS invPEs_1_3 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_1_3_io_in),
    .io_out(invPEs_1_3_io_out)
  );
  AES_InvS invPEs_2_0 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_2_0_io_in),
    .io_out(invPEs_2_0_io_out)
  );
  AES_InvS invPEs_2_1 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_2_1_io_in),
    .io_out(invPEs_2_1_io_out)
  );
  AES_InvS invPEs_2_2 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_2_2_io_in),
    .io_out(invPEs_2_2_io_out)
  );
  AES_InvS invPEs_2_3 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_2_3_io_in),
    .io_out(invPEs_2_3_io_out)
  );
  AES_InvS invPEs_3_0 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_3_0_io_in),
    .io_out(invPEs_3_0_io_out)
  );
  AES_InvS invPEs_3_1 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_3_1_io_in),
    .io_out(invPEs_3_1_io_out)
  );
  AES_InvS invPEs_3_2 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_3_2_io_in),
    .io_out(invPEs_3_2_io_out)
  );
  AES_InvS invPEs_3_3 ( // @[AES_PipelinedElasticBuffer.scala 689:22]
    .io_in(invPEs_3_3_io_in),
    .io_out(invPEs_3_3_io_out)
  );
  assign io_out_state_0_0 = invPEs_0_0_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_0_1 = invPEs_0_1_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_0_2 = invPEs_0_2_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_0_3 = invPEs_0_3_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_1_0 = invPEs_1_0_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_1_1 = invPEs_1_1_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_1_2 = invPEs_1_2_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_1_3 = invPEs_1_3_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_2_0 = invPEs_2_0_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_2_1 = invPEs_2_1_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_2_2 = invPEs_2_2_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_2_3 = invPEs_2_3_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_3_0 = invPEs_3_0_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_3_1 = invPEs_3_1_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_3_2 = invPEs_3_2_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign io_out_state_3_3 = invPEs_3_3_io_out; // @[AES_PipelinedElasticBuffer.scala 698:28]
  assign invPEs_0_0_io_in = io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_0_1_io_in = io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_0_2_io_in = io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_0_3_io_in = io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_1_0_io_in = io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_1_1_io_in = io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_1_2_io_in = io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_1_3_io_in = io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_2_0_io_in = io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_2_1_io_in = io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_2_2_io_in = io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_2_3_io_in = io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_3_0_io_in = io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_3_1_io_in = io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_3_2_io_in = io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 697:28]
  assign invPEs_3_3_io_in = io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 697:28]
endmodule
module AES_RotWord(
  output [31:0] io_out,
  input  [31:0] io_in
);
  wire [23:0] hi = io_in[23:0]; // @[AES_PipelinedElasticBuffer.scala 356:22]
  wire [7:0] lo = io_in[31:24]; // @[AES_PipelinedElasticBuffer.scala 356:35]
  assign io_out = {hi,lo}; // @[Cat.scala 30:58]
endmodule
module AES_SubWord(
  output [31:0] io_out,
  input  [31:0] io_in
);
  wire [7:0] PEs_0_io_in; // @[AES_PipelinedElasticBuffer.scala 342:20]
  wire [7:0] PEs_0_io_out; // @[AES_PipelinedElasticBuffer.scala 342:20]
  wire [7:0] PEs_1_io_in; // @[AES_PipelinedElasticBuffer.scala 342:20]
  wire [7:0] PEs_1_io_out; // @[AES_PipelinedElasticBuffer.scala 342:20]
  wire [7:0] PEs_2_io_in; // @[AES_PipelinedElasticBuffer.scala 342:20]
  wire [7:0] PEs_2_io_out; // @[AES_PipelinedElasticBuffer.scala 342:20]
  wire [7:0] PEs_3_io_in; // @[AES_PipelinedElasticBuffer.scala 342:20]
  wire [7:0] PEs_3_io_out; // @[AES_PipelinedElasticBuffer.scala 342:20]
  wire [15:0] lo = {PEs_1_io_out,PEs_0_io_out}; // @[Cat.scala 30:58]
  wire [15:0] hi = {PEs_3_io_out,PEs_2_io_out}; // @[Cat.scala 30:58]
  AES_S PEs_0 ( // @[AES_PipelinedElasticBuffer.scala 342:20]
    .io_in(PEs_0_io_in),
    .io_out(PEs_0_io_out)
  );
  AES_S PEs_1 ( // @[AES_PipelinedElasticBuffer.scala 342:20]
    .io_in(PEs_1_io_in),
    .io_out(PEs_1_io_out)
  );
  AES_S PEs_2 ( // @[AES_PipelinedElasticBuffer.scala 342:20]
    .io_in(PEs_2_io_in),
    .io_out(PEs_2_io_out)
  );
  AES_S PEs_3 ( // @[AES_PipelinedElasticBuffer.scala 342:20]
    .io_in(PEs_3_io_in),
    .io_out(PEs_3_io_out)
  );
  assign io_out = {hi,lo}; // @[Cat.scala 30:58]
  assign PEs_0_io_in = io_in[7:0]; // @[AES_PipelinedElasticBuffer.scala 343:22]
  assign PEs_1_io_in = io_in[15:8]; // @[AES_PipelinedElasticBuffer.scala 343:22]
  assign PEs_2_io_in = io_in[23:16]; // @[AES_PipelinedElasticBuffer.scala 343:22]
  assign PEs_3_io_in = io_in[31:24]; // @[AES_PipelinedElasticBuffer.scala 343:22]
endmodule
module AES_GetNewKey(
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 237:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 240:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 241:13]
endmodule
module AES_InvGetNewKey(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] w4 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w5 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w6 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [31:0] w7 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] w3 = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  wire [31:0] w2 = w6 ^ w5; // @[AES_PipelinedElasticBuffer.scala 301:12]
  wire [31:0] w1 = w5 ^ w4; // @[AES_PipelinedElasticBuffer.scala 302:12]
  wire [31:0] temp = 32'h36000000 ^ sub_io_out; // @[AES_PipelinedElasticBuffer.scala 310:16]
  wire [31:0] w0 = w4 ^ temp; // @[AES_PipelinedElasticBuffer.scala 303:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 305:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 308:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w0[31:24]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_1 = w0[23:16]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_2 = w0[15:8]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_3 = w0[7:0]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_1_0 = w1[31:24]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_1 = w1[23:16]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_2 = w1[15:8]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_3 = w1[7:0]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_2_0 = w2[31:24]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_1 = w2[23:16]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_2 = w2[15:8]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_3 = w2[7:0]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_3_0 = w3[31:24]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_1 = w3[23:16]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_2 = w3[15:8]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_3 = w3[7:0]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign rot_io_in = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 309:13]
endmodule
module AES_ProcessingElement(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 146:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:23 AES_PipelinedElasticBuffer.scala 156:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 163:21 AES_PipelinedElasticBuffer.scala 163:21]
  AES_XOR xor_ ( // @[AES_PipelinedElasticBuffer.scala 169:19]
    .io_out_state_0_0(xor__io_out_state_0_0),
    .io_out_state_0_1(xor__io_out_state_0_1),
    .io_out_state_0_2(xor__io_out_state_0_2),
    .io_out_state_0_3(xor__io_out_state_0_3),
    .io_out_state_1_0(xor__io_out_state_1_0),
    .io_out_state_1_1(xor__io_out_state_1_1),
    .io_out_state_1_2(xor__io_out_state_1_2),
    .io_out_state_1_3(xor__io_out_state_1_3),
    .io_out_state_2_0(xor__io_out_state_2_0),
    .io_out_state_2_1(xor__io_out_state_2_1),
    .io_out_state_2_2(xor__io_out_state_2_2),
    .io_out_state_2_3(xor__io_out_state_2_3),
    .io_out_state_3_0(xor__io_out_state_3_0),
    .io_out_state_3_1(xor__io_out_state_3_1),
    .io_out_state_3_2(xor__io_out_state_3_2),
    .io_out_state_3_3(xor__io_out_state_3_3),
    .io_in_state_0_0(xor__io_in_state_0_0),
    .io_in_state_0_1(xor__io_in_state_0_1),
    .io_in_state_0_2(xor__io_in_state_0_2),
    .io_in_state_0_3(xor__io_in_state_0_3),
    .io_in_state_1_0(xor__io_in_state_1_0),
    .io_in_state_1_1(xor__io_in_state_1_1),
    .io_in_state_1_2(xor__io_in_state_1_2),
    .io_in_state_1_3(xor__io_in_state_1_3),
    .io_in_state_2_0(xor__io_in_state_2_0),
    .io_in_state_2_1(xor__io_in_state_2_1),
    .io_in_state_2_2(xor__io_in_state_2_2),
    .io_in_state_2_3(xor__io_in_state_2_3),
    .io_in_state_3_0(xor__io_in_state_3_0),
    .io_in_state_3_1(xor__io_in_state_3_1),
    .io_in_state_3_2(xor__io_in_state_3_2),
    .io_in_state_3_3(xor__io_in_state_3_3),
    .io_in_key_0_0(xor__io_in_key_0_0),
    .io_in_key_0_1(xor__io_in_key_0_1),
    .io_in_key_0_2(xor__io_in_key_0_2),
    .io_in_key_0_3(xor__io_in_key_0_3),
    .io_in_key_1_0(xor__io_in_key_1_0),
    .io_in_key_1_1(xor__io_in_key_1_1),
    .io_in_key_1_2(xor__io_in_key_1_2),
    .io_in_key_1_3(xor__io_in_key_1_3),
    .io_in_key_2_0(xor__io_in_key_2_0),
    .io_in_key_2_1(xor__io_in_key_2_1),
    .io_in_key_2_2(xor__io_in_key_2_2),
    .io_in_key_2_3(xor__io_in_key_2_3),
    .io_in_key_3_0(xor__io_in_key_3_0),
    .io_in_key_3_1(xor__io_in_key_3_1),
    .io_in_key_3_2(xor__io_in_key_3_2),
    .io_in_key_3_3(xor__io_in_key_3_3)
  );
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 174:19]
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_XOR invxor ( // @[AES_PipelinedElasticBuffer.scala 184:22]
    .io_out_state_0_0(invxor_io_out_state_0_0),
    .io_out_state_0_1(invxor_io_out_state_0_1),
    .io_out_state_0_2(invxor_io_out_state_0_2),
    .io_out_state_0_3(invxor_io_out_state_0_3),
    .io_out_state_1_0(invxor_io_out_state_1_0),
    .io_out_state_1_1(invxor_io_out_state_1_1),
    .io_out_state_1_2(invxor_io_out_state_1_2),
    .io_out_state_1_3(invxor_io_out_state_1_3),
    .io_out_state_2_0(invxor_io_out_state_2_0),
    .io_out_state_2_1(invxor_io_out_state_2_1),
    .io_out_state_2_2(invxor_io_out_state_2_2),
    .io_out_state_2_3(invxor_io_out_state_2_3),
    .io_out_state_3_0(invxor_io_out_state_3_0),
    .io_out_state_3_1(invxor_io_out_state_3_1),
    .io_out_state_3_2(invxor_io_out_state_3_2),
    .io_out_state_3_3(invxor_io_out_state_3_3),
    .io_in_state_0_0(invxor_io_in_state_0_0),
    .io_in_state_0_1(invxor_io_in_state_0_1),
    .io_in_state_0_2(invxor_io_in_state_0_2),
    .io_in_state_0_3(invxor_io_in_state_0_3),
    .io_in_state_1_0(invxor_io_in_state_1_0),
    .io_in_state_1_1(invxor_io_in_state_1_1),
    .io_in_state_1_2(invxor_io_in_state_1_2),
    .io_in_state_1_3(invxor_io_in_state_1_3),
    .io_in_state_2_0(invxor_io_in_state_2_0),
    .io_in_state_2_1(invxor_io_in_state_2_1),
    .io_in_state_2_2(invxor_io_in_state_2_2),
    .io_in_state_2_3(invxor_io_in_state_2_3),
    .io_in_state_3_0(invxor_io_in_state_3_0),
    .io_in_state_3_1(invxor_io_in_state_3_1),
    .io_in_state_3_2(invxor_io_in_state_3_2),
    .io_in_state_3_3(invxor_io_in_state_3_3),
    .io_in_key_0_0(invxor_io_in_key_0_0),
    .io_in_key_0_1(invxor_io_in_key_0_1),
    .io_in_key_0_2(invxor_io_in_key_0_2),
    .io_in_key_0_3(invxor_io_in_key_0_3),
    .io_in_key_1_0(invxor_io_in_key_1_0),
    .io_in_key_1_1(invxor_io_in_key_1_1),
    .io_in_key_1_2(invxor_io_in_key_1_2),
    .io_in_key_1_3(invxor_io_in_key_1_3),
    .io_in_key_2_0(invxor_io_in_key_2_0),
    .io_in_key_2_1(invxor_io_in_key_2_1),
    .io_in_key_2_2(invxor_io_in_key_2_2),
    .io_in_key_2_3(invxor_io_in_key_2_3),
    .io_in_key_3_0(invxor_io_in_key_3_0),
    .io_in_key_3_1(invxor_io_in_key_3_1),
    .io_in_key_3_2(invxor_io_in_key_3_2),
    .io_in_key_3_3(invxor_io_in_key_3_3)
  );
  AES_InvMixColumns invmix ( // @[AES_PipelinedElasticBuffer.scala 189:22]
    .io_out_state_0_0(invmix_io_out_state_0_0),
    .io_out_state_0_1(invmix_io_out_state_0_1),
    .io_out_state_0_2(invmix_io_out_state_0_2),
    .io_out_state_0_3(invmix_io_out_state_0_3),
    .io_out_state_1_0(invmix_io_out_state_1_0),
    .io_out_state_1_1(invmix_io_out_state_1_1),
    .io_out_state_1_2(invmix_io_out_state_1_2),
    .io_out_state_1_3(invmix_io_out_state_1_3),
    .io_out_state_2_0(invmix_io_out_state_2_0),
    .io_out_state_2_1(invmix_io_out_state_2_1),
    .io_out_state_2_2(invmix_io_out_state_2_2),
    .io_out_state_2_3(invmix_io_out_state_2_3),
    .io_out_state_3_0(invmix_io_out_state_3_0),
    .io_out_state_3_1(invmix_io_out_state_3_1),
    .io_out_state_3_2(invmix_io_out_state_3_2),
    .io_out_state_3_3(invmix_io_out_state_3_3),
    .io_in_state_0_0(invmix_io_in_state_0_0),
    .io_in_state_0_1(invmix_io_in_state_0_1),
    .io_in_state_0_2(invmix_io_in_state_0_2),
    .io_in_state_0_3(invmix_io_in_state_0_3),
    .io_in_state_1_0(invmix_io_in_state_1_0),
    .io_in_state_1_1(invmix_io_in_state_1_1),
    .io_in_state_1_2(invmix_io_in_state_1_2),
    .io_in_state_1_3(invmix_io_in_state_1_3),
    .io_in_state_2_0(invmix_io_in_state_2_0),
    .io_in_state_2_1(invmix_io_in_state_2_1),
    .io_in_state_2_2(invmix_io_in_state_2_2),
    .io_in_state_2_3(invmix_io_in_state_2_3),
    .io_in_state_3_0(invmix_io_in_state_3_0),
    .io_in_state_3_1(invmix_io_in_state_3_1),
    .io_in_state_3_2(invmix_io_in_state_3_2),
    .io_in_state_3_3(invmix_io_in_state_3_3)
  );
  AES_InvShiftRows invshift ( // @[AES_PipelinedElasticBuffer.scala 192:24]
    .io_out_state_0_0(invshift_io_out_state_0_0),
    .io_out_state_0_1(invshift_io_out_state_0_1),
    .io_out_state_0_2(invshift_io_out_state_0_2),
    .io_out_state_0_3(invshift_io_out_state_0_3),
    .io_out_state_1_0(invshift_io_out_state_1_0),
    .io_out_state_1_1(invshift_io_out_state_1_1),
    .io_out_state_1_2(invshift_io_out_state_1_2),
    .io_out_state_1_3(invshift_io_out_state_1_3),
    .io_out_state_2_0(invshift_io_out_state_2_0),
    .io_out_state_2_1(invshift_io_out_state_2_1),
    .io_out_state_2_2(invshift_io_out_state_2_2),
    .io_out_state_2_3(invshift_io_out_state_2_3),
    .io_out_state_3_0(invshift_io_out_state_3_0),
    .io_out_state_3_1(invshift_io_out_state_3_1),
    .io_out_state_3_2(invshift_io_out_state_3_2),
    .io_out_state_3_3(invshift_io_out_state_3_3),
    .io_in_state_0_0(invshift_io_in_state_0_0),
    .io_in_state_0_1(invshift_io_in_state_0_1),
    .io_in_state_0_2(invshift_io_in_state_0_2),
    .io_in_state_0_3(invshift_io_in_state_0_3),
    .io_in_state_1_0(invshift_io_in_state_1_0),
    .io_in_state_1_1(invshift_io_in_state_1_1),
    .io_in_state_1_2(invshift_io_in_state_1_2),
    .io_in_state_1_3(invshift_io_in_state_1_3),
    .io_in_state_2_0(invshift_io_in_state_2_0),
    .io_in_state_2_1(invshift_io_in_state_2_1),
    .io_in_state_2_2(invshift_io_in_state_2_2),
    .io_in_state_2_3(invshift_io_in_state_2_3),
    .io_in_state_3_0(invshift_io_in_state_3_0),
    .io_in_state_3_1(invshift_io_in_state_3_1),
    .io_in_state_3_2(invshift_io_in_state_3_2),
    .io_in_state_3_3(invshift_io_in_state_3_3)
  );
  AES_InvSubBytes invsub ( // @[AES_PipelinedElasticBuffer.scala 199:22]
    .io_out_state_0_0(invsub_io_out_state_0_0),
    .io_out_state_0_1(invsub_io_out_state_0_1),
    .io_out_state_0_2(invsub_io_out_state_0_2),
    .io_out_state_0_3(invsub_io_out_state_0_3),
    .io_out_state_1_0(invsub_io_out_state_1_0),
    .io_out_state_1_1(invsub_io_out_state_1_1),
    .io_out_state_1_2(invsub_io_out_state_1_2),
    .io_out_state_1_3(invsub_io_out_state_1_3),
    .io_out_state_2_0(invsub_io_out_state_2_0),
    .io_out_state_2_1(invsub_io_out_state_2_1),
    .io_out_state_2_2(invsub_io_out_state_2_2),
    .io_out_state_2_3(invsub_io_out_state_2_3),
    .io_out_state_3_0(invsub_io_out_state_3_0),
    .io_out_state_3_1(invsub_io_out_state_3_1),
    .io_out_state_3_2(invsub_io_out_state_3_2),
    .io_out_state_3_3(invsub_io_out_state_3_3),
    .io_in_state_0_0(invsub_io_in_state_0_0),
    .io_in_state_0_1(invsub_io_in_state_0_1),
    .io_in_state_0_2(invsub_io_in_state_0_2),
    .io_in_state_0_3(invsub_io_in_state_0_3),
    .io_in_state_1_0(invsub_io_in_state_1_0),
    .io_in_state_1_1(invsub_io_in_state_1_1),
    .io_in_state_1_2(invsub_io_in_state_1_2),
    .io_in_state_1_3(invsub_io_in_state_1_3),
    .io_in_state_2_0(invsub_io_in_state_2_0),
    .io_in_state_2_1(invsub_io_in_state_2_1),
    .io_in_state_2_2(invsub_io_in_state_2_2),
    .io_in_state_2_3(invsub_io_in_state_2_3),
    .io_in_state_3_0(invsub_io_in_state_3_0),
    .io_in_state_3_1(invsub_io_in_state_3_1),
    .io_in_state_3_2(invsub_io_in_state_3_2),
    .io_in_state_3_3(invsub_io_in_state_3_3)
  );
  AES_GetNewKey key ( // @[AES_PipelinedElasticBuffer.scala 202:19]
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  AES_InvGetNewKey invkey ( // @[AES_PipelinedElasticBuffer.scala 206:22]
    .io_out_key_0_0(invkey_io_out_key_0_0),
    .io_out_key_0_1(invkey_io_out_key_0_1),
    .io_out_key_0_2(invkey_io_out_key_0_2),
    .io_out_key_0_3(invkey_io_out_key_0_3),
    .io_out_key_1_0(invkey_io_out_key_1_0),
    .io_out_key_1_1(invkey_io_out_key_1_1),
    .io_out_key_1_2(invkey_io_out_key_1_2),
    .io_out_key_1_3(invkey_io_out_key_1_3),
    .io_out_key_2_0(invkey_io_out_key_2_0),
    .io_out_key_2_1(invkey_io_out_key_2_1),
    .io_out_key_2_2(invkey_io_out_key_2_2),
    .io_out_key_2_3(invkey_io_out_key_2_3),
    .io_out_key_3_0(invkey_io_out_key_3_0),
    .io_out_key_3_1(invkey_io_out_key_3_1),
    .io_out_key_3_2(invkey_io_out_key_3_2),
    .io_out_key_3_3(invkey_io_out_key_3_3),
    .io_in_key_0_0(invkey_io_in_key_0_0),
    .io_in_key_0_1(invkey_io_in_key_0_1),
    .io_in_key_0_2(invkey_io_in_key_0_2),
    .io_in_key_0_3(invkey_io_in_key_0_3),
    .io_in_key_1_0(invkey_io_in_key_1_0),
    .io_in_key_1_1(invkey_io_in_key_1_1),
    .io_in_key_1_2(invkey_io_in_key_1_2),
    .io_in_key_1_3(invkey_io_in_key_1_3),
    .io_in_key_2_0(invkey_io_in_key_2_0),
    .io_in_key_2_1(invkey_io_in_key_2_1),
    .io_in_key_2_2(invkey_io_in_key_2_2),
    .io_in_key_2_3(invkey_io_in_key_2_3),
    .io_in_key_3_0(invkey_io_in_key_3_0),
    .io_in_key_3_1(invkey_io_in_key_3_1),
    .io_in_key_3_2(invkey_io_in_key_3_2),
    .io_in_key_3_3(invkey_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 151:27]
  assign io_out_bits_state_0_0 = invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_1 = invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_2 = invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_3 = invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_0 = invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_1 = invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_2 = invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_3 = invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_0 = invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_1 = invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_2 = invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_3 = invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_0 = invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_1 = invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_2 = invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_3 = invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_0 = invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_1 = invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_2 = invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_3 = invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_0 = invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_1 = invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_2 = invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_3 = invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_0 = invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_1 = invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_2 = invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_3 = invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_0 = invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_1 = invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_2 = invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_3 = invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 150:18]
  assign xor__io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign sub_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign invxor_io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invmix_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invshift_io_in_state_0_0 = invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_0_1 = invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_0_2 = invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_0_3 = invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_1_0 = invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_1_1 = invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_1_2 = invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_1_3 = invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_2_0 = invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_2_1 = invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_2_2 = invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_2_3 = invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_3_0 = invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_3_1 = invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_3_2 = invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invshift_io_in_state_3_3 = invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 194:20]
  assign invsub_io_in_state_0_0 = invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_1 = invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_2 = invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_3 = invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_0 = invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_1 = invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_2 = invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_3 = invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_0 = invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_1 = invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_2 = invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_3 = invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_0 = invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_1 = invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_2 = invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_3 = invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 146:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 146:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 165:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 159:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_1(
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 237:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 240:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 241:13]
endmodule
module AES_InvGetNewKey_1(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] w4 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w5 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w6 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [31:0] w7 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] w3 = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  wire [31:0] w2 = w6 ^ w5; // @[AES_PipelinedElasticBuffer.scala 301:12]
  wire [31:0] w1 = w5 ^ w4; // @[AES_PipelinedElasticBuffer.scala 302:12]
  wire [31:0] temp = 32'h1b000000 ^ sub_io_out; // @[AES_PipelinedElasticBuffer.scala 310:16]
  wire [31:0] w0 = w4 ^ temp; // @[AES_PipelinedElasticBuffer.scala 303:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 305:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 308:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w0[31:24]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_1 = w0[23:16]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_2 = w0[15:8]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_3 = w0[7:0]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_1_0 = w1[31:24]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_1 = w1[23:16]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_2 = w1[15:8]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_3 = w1[7:0]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_2_0 = w2[31:24]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_1 = w2[23:16]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_2 = w2[15:8]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_3 = w2[7:0]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_3_0 = w3[31:24]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_1 = w3[23:16]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_2 = w3[15:8]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_3 = w3[7:0]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign rot_io_in = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 309:13]
endmodule
module AES_ProcessingElement_1(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 146:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:23 AES_PipelinedElasticBuffer.scala 156:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 163:21 AES_PipelinedElasticBuffer.scala 163:21]
  AES_XOR xor_ ( // @[AES_PipelinedElasticBuffer.scala 169:19]
    .io_out_state_0_0(xor__io_out_state_0_0),
    .io_out_state_0_1(xor__io_out_state_0_1),
    .io_out_state_0_2(xor__io_out_state_0_2),
    .io_out_state_0_3(xor__io_out_state_0_3),
    .io_out_state_1_0(xor__io_out_state_1_0),
    .io_out_state_1_1(xor__io_out_state_1_1),
    .io_out_state_1_2(xor__io_out_state_1_2),
    .io_out_state_1_3(xor__io_out_state_1_3),
    .io_out_state_2_0(xor__io_out_state_2_0),
    .io_out_state_2_1(xor__io_out_state_2_1),
    .io_out_state_2_2(xor__io_out_state_2_2),
    .io_out_state_2_3(xor__io_out_state_2_3),
    .io_out_state_3_0(xor__io_out_state_3_0),
    .io_out_state_3_1(xor__io_out_state_3_1),
    .io_out_state_3_2(xor__io_out_state_3_2),
    .io_out_state_3_3(xor__io_out_state_3_3),
    .io_in_state_0_0(xor__io_in_state_0_0),
    .io_in_state_0_1(xor__io_in_state_0_1),
    .io_in_state_0_2(xor__io_in_state_0_2),
    .io_in_state_0_3(xor__io_in_state_0_3),
    .io_in_state_1_0(xor__io_in_state_1_0),
    .io_in_state_1_1(xor__io_in_state_1_1),
    .io_in_state_1_2(xor__io_in_state_1_2),
    .io_in_state_1_3(xor__io_in_state_1_3),
    .io_in_state_2_0(xor__io_in_state_2_0),
    .io_in_state_2_1(xor__io_in_state_2_1),
    .io_in_state_2_2(xor__io_in_state_2_2),
    .io_in_state_2_3(xor__io_in_state_2_3),
    .io_in_state_3_0(xor__io_in_state_3_0),
    .io_in_state_3_1(xor__io_in_state_3_1),
    .io_in_state_3_2(xor__io_in_state_3_2),
    .io_in_state_3_3(xor__io_in_state_3_3),
    .io_in_key_0_0(xor__io_in_key_0_0),
    .io_in_key_0_1(xor__io_in_key_0_1),
    .io_in_key_0_2(xor__io_in_key_0_2),
    .io_in_key_0_3(xor__io_in_key_0_3),
    .io_in_key_1_0(xor__io_in_key_1_0),
    .io_in_key_1_1(xor__io_in_key_1_1),
    .io_in_key_1_2(xor__io_in_key_1_2),
    .io_in_key_1_3(xor__io_in_key_1_3),
    .io_in_key_2_0(xor__io_in_key_2_0),
    .io_in_key_2_1(xor__io_in_key_2_1),
    .io_in_key_2_2(xor__io_in_key_2_2),
    .io_in_key_2_3(xor__io_in_key_2_3),
    .io_in_key_3_0(xor__io_in_key_3_0),
    .io_in_key_3_1(xor__io_in_key_3_1),
    .io_in_key_3_2(xor__io_in_key_3_2),
    .io_in_key_3_3(xor__io_in_key_3_3)
  );
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 174:19]
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_XOR invxor ( // @[AES_PipelinedElasticBuffer.scala 184:22]
    .io_out_state_0_0(invxor_io_out_state_0_0),
    .io_out_state_0_1(invxor_io_out_state_0_1),
    .io_out_state_0_2(invxor_io_out_state_0_2),
    .io_out_state_0_3(invxor_io_out_state_0_3),
    .io_out_state_1_0(invxor_io_out_state_1_0),
    .io_out_state_1_1(invxor_io_out_state_1_1),
    .io_out_state_1_2(invxor_io_out_state_1_2),
    .io_out_state_1_3(invxor_io_out_state_1_3),
    .io_out_state_2_0(invxor_io_out_state_2_0),
    .io_out_state_2_1(invxor_io_out_state_2_1),
    .io_out_state_2_2(invxor_io_out_state_2_2),
    .io_out_state_2_3(invxor_io_out_state_2_3),
    .io_out_state_3_0(invxor_io_out_state_3_0),
    .io_out_state_3_1(invxor_io_out_state_3_1),
    .io_out_state_3_2(invxor_io_out_state_3_2),
    .io_out_state_3_3(invxor_io_out_state_3_3),
    .io_in_state_0_0(invxor_io_in_state_0_0),
    .io_in_state_0_1(invxor_io_in_state_0_1),
    .io_in_state_0_2(invxor_io_in_state_0_2),
    .io_in_state_0_3(invxor_io_in_state_0_3),
    .io_in_state_1_0(invxor_io_in_state_1_0),
    .io_in_state_1_1(invxor_io_in_state_1_1),
    .io_in_state_1_2(invxor_io_in_state_1_2),
    .io_in_state_1_3(invxor_io_in_state_1_3),
    .io_in_state_2_0(invxor_io_in_state_2_0),
    .io_in_state_2_1(invxor_io_in_state_2_1),
    .io_in_state_2_2(invxor_io_in_state_2_2),
    .io_in_state_2_3(invxor_io_in_state_2_3),
    .io_in_state_3_0(invxor_io_in_state_3_0),
    .io_in_state_3_1(invxor_io_in_state_3_1),
    .io_in_state_3_2(invxor_io_in_state_3_2),
    .io_in_state_3_3(invxor_io_in_state_3_3),
    .io_in_key_0_0(invxor_io_in_key_0_0),
    .io_in_key_0_1(invxor_io_in_key_0_1),
    .io_in_key_0_2(invxor_io_in_key_0_2),
    .io_in_key_0_3(invxor_io_in_key_0_3),
    .io_in_key_1_0(invxor_io_in_key_1_0),
    .io_in_key_1_1(invxor_io_in_key_1_1),
    .io_in_key_1_2(invxor_io_in_key_1_2),
    .io_in_key_1_3(invxor_io_in_key_1_3),
    .io_in_key_2_0(invxor_io_in_key_2_0),
    .io_in_key_2_1(invxor_io_in_key_2_1),
    .io_in_key_2_2(invxor_io_in_key_2_2),
    .io_in_key_2_3(invxor_io_in_key_2_3),
    .io_in_key_3_0(invxor_io_in_key_3_0),
    .io_in_key_3_1(invxor_io_in_key_3_1),
    .io_in_key_3_2(invxor_io_in_key_3_2),
    .io_in_key_3_3(invxor_io_in_key_3_3)
  );
  AES_InvMixColumns invmix ( // @[AES_PipelinedElasticBuffer.scala 189:22]
    .io_out_state_0_0(invmix_io_out_state_0_0),
    .io_out_state_0_1(invmix_io_out_state_0_1),
    .io_out_state_0_2(invmix_io_out_state_0_2),
    .io_out_state_0_3(invmix_io_out_state_0_3),
    .io_out_state_1_0(invmix_io_out_state_1_0),
    .io_out_state_1_1(invmix_io_out_state_1_1),
    .io_out_state_1_2(invmix_io_out_state_1_2),
    .io_out_state_1_3(invmix_io_out_state_1_3),
    .io_out_state_2_0(invmix_io_out_state_2_0),
    .io_out_state_2_1(invmix_io_out_state_2_1),
    .io_out_state_2_2(invmix_io_out_state_2_2),
    .io_out_state_2_3(invmix_io_out_state_2_3),
    .io_out_state_3_0(invmix_io_out_state_3_0),
    .io_out_state_3_1(invmix_io_out_state_3_1),
    .io_out_state_3_2(invmix_io_out_state_3_2),
    .io_out_state_3_3(invmix_io_out_state_3_3),
    .io_in_state_0_0(invmix_io_in_state_0_0),
    .io_in_state_0_1(invmix_io_in_state_0_1),
    .io_in_state_0_2(invmix_io_in_state_0_2),
    .io_in_state_0_3(invmix_io_in_state_0_3),
    .io_in_state_1_0(invmix_io_in_state_1_0),
    .io_in_state_1_1(invmix_io_in_state_1_1),
    .io_in_state_1_2(invmix_io_in_state_1_2),
    .io_in_state_1_3(invmix_io_in_state_1_3),
    .io_in_state_2_0(invmix_io_in_state_2_0),
    .io_in_state_2_1(invmix_io_in_state_2_1),
    .io_in_state_2_2(invmix_io_in_state_2_2),
    .io_in_state_2_3(invmix_io_in_state_2_3),
    .io_in_state_3_0(invmix_io_in_state_3_0),
    .io_in_state_3_1(invmix_io_in_state_3_1),
    .io_in_state_3_2(invmix_io_in_state_3_2),
    .io_in_state_3_3(invmix_io_in_state_3_3)
  );
  AES_InvShiftRows invshift ( // @[AES_PipelinedElasticBuffer.scala 192:24]
    .io_out_state_0_0(invshift_io_out_state_0_0),
    .io_out_state_0_1(invshift_io_out_state_0_1),
    .io_out_state_0_2(invshift_io_out_state_0_2),
    .io_out_state_0_3(invshift_io_out_state_0_3),
    .io_out_state_1_0(invshift_io_out_state_1_0),
    .io_out_state_1_1(invshift_io_out_state_1_1),
    .io_out_state_1_2(invshift_io_out_state_1_2),
    .io_out_state_1_3(invshift_io_out_state_1_3),
    .io_out_state_2_0(invshift_io_out_state_2_0),
    .io_out_state_2_1(invshift_io_out_state_2_1),
    .io_out_state_2_2(invshift_io_out_state_2_2),
    .io_out_state_2_3(invshift_io_out_state_2_3),
    .io_out_state_3_0(invshift_io_out_state_3_0),
    .io_out_state_3_1(invshift_io_out_state_3_1),
    .io_out_state_3_2(invshift_io_out_state_3_2),
    .io_out_state_3_3(invshift_io_out_state_3_3),
    .io_in_state_0_0(invshift_io_in_state_0_0),
    .io_in_state_0_1(invshift_io_in_state_0_1),
    .io_in_state_0_2(invshift_io_in_state_0_2),
    .io_in_state_0_3(invshift_io_in_state_0_3),
    .io_in_state_1_0(invshift_io_in_state_1_0),
    .io_in_state_1_1(invshift_io_in_state_1_1),
    .io_in_state_1_2(invshift_io_in_state_1_2),
    .io_in_state_1_3(invshift_io_in_state_1_3),
    .io_in_state_2_0(invshift_io_in_state_2_0),
    .io_in_state_2_1(invshift_io_in_state_2_1),
    .io_in_state_2_2(invshift_io_in_state_2_2),
    .io_in_state_2_3(invshift_io_in_state_2_3),
    .io_in_state_3_0(invshift_io_in_state_3_0),
    .io_in_state_3_1(invshift_io_in_state_3_1),
    .io_in_state_3_2(invshift_io_in_state_3_2),
    .io_in_state_3_3(invshift_io_in_state_3_3)
  );
  AES_InvSubBytes invsub ( // @[AES_PipelinedElasticBuffer.scala 199:22]
    .io_out_state_0_0(invsub_io_out_state_0_0),
    .io_out_state_0_1(invsub_io_out_state_0_1),
    .io_out_state_0_2(invsub_io_out_state_0_2),
    .io_out_state_0_3(invsub_io_out_state_0_3),
    .io_out_state_1_0(invsub_io_out_state_1_0),
    .io_out_state_1_1(invsub_io_out_state_1_1),
    .io_out_state_1_2(invsub_io_out_state_1_2),
    .io_out_state_1_3(invsub_io_out_state_1_3),
    .io_out_state_2_0(invsub_io_out_state_2_0),
    .io_out_state_2_1(invsub_io_out_state_2_1),
    .io_out_state_2_2(invsub_io_out_state_2_2),
    .io_out_state_2_3(invsub_io_out_state_2_3),
    .io_out_state_3_0(invsub_io_out_state_3_0),
    .io_out_state_3_1(invsub_io_out_state_3_1),
    .io_out_state_3_2(invsub_io_out_state_3_2),
    .io_out_state_3_3(invsub_io_out_state_3_3),
    .io_in_state_0_0(invsub_io_in_state_0_0),
    .io_in_state_0_1(invsub_io_in_state_0_1),
    .io_in_state_0_2(invsub_io_in_state_0_2),
    .io_in_state_0_3(invsub_io_in_state_0_3),
    .io_in_state_1_0(invsub_io_in_state_1_0),
    .io_in_state_1_1(invsub_io_in_state_1_1),
    .io_in_state_1_2(invsub_io_in_state_1_2),
    .io_in_state_1_3(invsub_io_in_state_1_3),
    .io_in_state_2_0(invsub_io_in_state_2_0),
    .io_in_state_2_1(invsub_io_in_state_2_1),
    .io_in_state_2_2(invsub_io_in_state_2_2),
    .io_in_state_2_3(invsub_io_in_state_2_3),
    .io_in_state_3_0(invsub_io_in_state_3_0),
    .io_in_state_3_1(invsub_io_in_state_3_1),
    .io_in_state_3_2(invsub_io_in_state_3_2),
    .io_in_state_3_3(invsub_io_in_state_3_3)
  );
  AES_GetNewKey_1 key ( // @[AES_PipelinedElasticBuffer.scala 202:19]
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  AES_InvGetNewKey_1 invkey ( // @[AES_PipelinedElasticBuffer.scala 206:22]
    .io_out_key_0_0(invkey_io_out_key_0_0),
    .io_out_key_0_1(invkey_io_out_key_0_1),
    .io_out_key_0_2(invkey_io_out_key_0_2),
    .io_out_key_0_3(invkey_io_out_key_0_3),
    .io_out_key_1_0(invkey_io_out_key_1_0),
    .io_out_key_1_1(invkey_io_out_key_1_1),
    .io_out_key_1_2(invkey_io_out_key_1_2),
    .io_out_key_1_3(invkey_io_out_key_1_3),
    .io_out_key_2_0(invkey_io_out_key_2_0),
    .io_out_key_2_1(invkey_io_out_key_2_1),
    .io_out_key_2_2(invkey_io_out_key_2_2),
    .io_out_key_2_3(invkey_io_out_key_2_3),
    .io_out_key_3_0(invkey_io_out_key_3_0),
    .io_out_key_3_1(invkey_io_out_key_3_1),
    .io_out_key_3_2(invkey_io_out_key_3_2),
    .io_out_key_3_3(invkey_io_out_key_3_3),
    .io_in_key_0_0(invkey_io_in_key_0_0),
    .io_in_key_0_1(invkey_io_in_key_0_1),
    .io_in_key_0_2(invkey_io_in_key_0_2),
    .io_in_key_0_3(invkey_io_in_key_0_3),
    .io_in_key_1_0(invkey_io_in_key_1_0),
    .io_in_key_1_1(invkey_io_in_key_1_1),
    .io_in_key_1_2(invkey_io_in_key_1_2),
    .io_in_key_1_3(invkey_io_in_key_1_3),
    .io_in_key_2_0(invkey_io_in_key_2_0),
    .io_in_key_2_1(invkey_io_in_key_2_1),
    .io_in_key_2_2(invkey_io_in_key_2_2),
    .io_in_key_2_3(invkey_io_in_key_2_3),
    .io_in_key_3_0(invkey_io_in_key_3_0),
    .io_in_key_3_1(invkey_io_in_key_3_1),
    .io_in_key_3_2(invkey_io_in_key_3_2),
    .io_in_key_3_3(invkey_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 151:27]
  assign io_out_bits_state_0_0 = invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_1 = invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_2 = invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_3 = invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_0 = invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_1 = invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_2 = invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_3 = invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_0 = invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_1 = invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_2 = invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_3 = invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_0 = invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_1 = invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_2 = invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_3 = invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_0 = invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_1 = invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_2 = invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_3 = invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_0 = invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_1 = invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_2 = invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_3 = invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_0 = invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_1 = invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_2 = invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_3 = invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_0 = invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_1 = invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_2 = invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_3 = invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 150:18]
  assign xor__io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign sub_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign invxor_io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invmix_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invshift_io_in_state_0_0 = invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_1 = invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_2 = invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_3 = invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_0 = invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_1 = invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_2 = invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_3 = invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_0 = invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_1 = invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_2 = invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_3 = invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_0 = invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_1 = invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_2 = invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_3 = invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invsub_io_in_state_0_0 = invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_1 = invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_2 = invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_3 = invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_0 = invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_1 = invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_2 = invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_3 = invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_0 = invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_1 = invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_2 = invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_3 = invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_0 = invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_1 = invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_2 = invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_3 = invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 146:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 146:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 165:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 159:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_2(
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 237:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 240:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 241:13]
endmodule
module AES_InvGetNewKey_2(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] w4 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w5 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w6 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [31:0] w7 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] w3 = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  wire [31:0] w2 = w6 ^ w5; // @[AES_PipelinedElasticBuffer.scala 301:12]
  wire [31:0] w1 = w5 ^ w4; // @[AES_PipelinedElasticBuffer.scala 302:12]
  wire [31:0] temp = 32'h80000000 ^ sub_io_out; // @[AES_PipelinedElasticBuffer.scala 310:16]
  wire [31:0] w0 = w4 ^ temp; // @[AES_PipelinedElasticBuffer.scala 303:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 305:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 308:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w0[31:24]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_1 = w0[23:16]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_2 = w0[15:8]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_3 = w0[7:0]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_1_0 = w1[31:24]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_1 = w1[23:16]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_2 = w1[15:8]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_3 = w1[7:0]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_2_0 = w2[31:24]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_1 = w2[23:16]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_2 = w2[15:8]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_3 = w2[7:0]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_3_0 = w3[31:24]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_1 = w3[23:16]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_2 = w3[15:8]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_3 = w3[7:0]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign rot_io_in = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 309:13]
endmodule
module AES_ProcessingElement_2(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 146:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:23 AES_PipelinedElasticBuffer.scala 156:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 163:21 AES_PipelinedElasticBuffer.scala 163:21]
  AES_XOR xor_ ( // @[AES_PipelinedElasticBuffer.scala 169:19]
    .io_out_state_0_0(xor__io_out_state_0_0),
    .io_out_state_0_1(xor__io_out_state_0_1),
    .io_out_state_0_2(xor__io_out_state_0_2),
    .io_out_state_0_3(xor__io_out_state_0_3),
    .io_out_state_1_0(xor__io_out_state_1_0),
    .io_out_state_1_1(xor__io_out_state_1_1),
    .io_out_state_1_2(xor__io_out_state_1_2),
    .io_out_state_1_3(xor__io_out_state_1_3),
    .io_out_state_2_0(xor__io_out_state_2_0),
    .io_out_state_2_1(xor__io_out_state_2_1),
    .io_out_state_2_2(xor__io_out_state_2_2),
    .io_out_state_2_3(xor__io_out_state_2_3),
    .io_out_state_3_0(xor__io_out_state_3_0),
    .io_out_state_3_1(xor__io_out_state_3_1),
    .io_out_state_3_2(xor__io_out_state_3_2),
    .io_out_state_3_3(xor__io_out_state_3_3),
    .io_in_state_0_0(xor__io_in_state_0_0),
    .io_in_state_0_1(xor__io_in_state_0_1),
    .io_in_state_0_2(xor__io_in_state_0_2),
    .io_in_state_0_3(xor__io_in_state_0_3),
    .io_in_state_1_0(xor__io_in_state_1_0),
    .io_in_state_1_1(xor__io_in_state_1_1),
    .io_in_state_1_2(xor__io_in_state_1_2),
    .io_in_state_1_3(xor__io_in_state_1_3),
    .io_in_state_2_0(xor__io_in_state_2_0),
    .io_in_state_2_1(xor__io_in_state_2_1),
    .io_in_state_2_2(xor__io_in_state_2_2),
    .io_in_state_2_3(xor__io_in_state_2_3),
    .io_in_state_3_0(xor__io_in_state_3_0),
    .io_in_state_3_1(xor__io_in_state_3_1),
    .io_in_state_3_2(xor__io_in_state_3_2),
    .io_in_state_3_3(xor__io_in_state_3_3),
    .io_in_key_0_0(xor__io_in_key_0_0),
    .io_in_key_0_1(xor__io_in_key_0_1),
    .io_in_key_0_2(xor__io_in_key_0_2),
    .io_in_key_0_3(xor__io_in_key_0_3),
    .io_in_key_1_0(xor__io_in_key_1_0),
    .io_in_key_1_1(xor__io_in_key_1_1),
    .io_in_key_1_2(xor__io_in_key_1_2),
    .io_in_key_1_3(xor__io_in_key_1_3),
    .io_in_key_2_0(xor__io_in_key_2_0),
    .io_in_key_2_1(xor__io_in_key_2_1),
    .io_in_key_2_2(xor__io_in_key_2_2),
    .io_in_key_2_3(xor__io_in_key_2_3),
    .io_in_key_3_0(xor__io_in_key_3_0),
    .io_in_key_3_1(xor__io_in_key_3_1),
    .io_in_key_3_2(xor__io_in_key_3_2),
    .io_in_key_3_3(xor__io_in_key_3_3)
  );
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 174:19]
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_XOR invxor ( // @[AES_PipelinedElasticBuffer.scala 184:22]
    .io_out_state_0_0(invxor_io_out_state_0_0),
    .io_out_state_0_1(invxor_io_out_state_0_1),
    .io_out_state_0_2(invxor_io_out_state_0_2),
    .io_out_state_0_3(invxor_io_out_state_0_3),
    .io_out_state_1_0(invxor_io_out_state_1_0),
    .io_out_state_1_1(invxor_io_out_state_1_1),
    .io_out_state_1_2(invxor_io_out_state_1_2),
    .io_out_state_1_3(invxor_io_out_state_1_3),
    .io_out_state_2_0(invxor_io_out_state_2_0),
    .io_out_state_2_1(invxor_io_out_state_2_1),
    .io_out_state_2_2(invxor_io_out_state_2_2),
    .io_out_state_2_3(invxor_io_out_state_2_3),
    .io_out_state_3_0(invxor_io_out_state_3_0),
    .io_out_state_3_1(invxor_io_out_state_3_1),
    .io_out_state_3_2(invxor_io_out_state_3_2),
    .io_out_state_3_3(invxor_io_out_state_3_3),
    .io_in_state_0_0(invxor_io_in_state_0_0),
    .io_in_state_0_1(invxor_io_in_state_0_1),
    .io_in_state_0_2(invxor_io_in_state_0_2),
    .io_in_state_0_3(invxor_io_in_state_0_3),
    .io_in_state_1_0(invxor_io_in_state_1_0),
    .io_in_state_1_1(invxor_io_in_state_1_1),
    .io_in_state_1_2(invxor_io_in_state_1_2),
    .io_in_state_1_3(invxor_io_in_state_1_3),
    .io_in_state_2_0(invxor_io_in_state_2_0),
    .io_in_state_2_1(invxor_io_in_state_2_1),
    .io_in_state_2_2(invxor_io_in_state_2_2),
    .io_in_state_2_3(invxor_io_in_state_2_3),
    .io_in_state_3_0(invxor_io_in_state_3_0),
    .io_in_state_3_1(invxor_io_in_state_3_1),
    .io_in_state_3_2(invxor_io_in_state_3_2),
    .io_in_state_3_3(invxor_io_in_state_3_3),
    .io_in_key_0_0(invxor_io_in_key_0_0),
    .io_in_key_0_1(invxor_io_in_key_0_1),
    .io_in_key_0_2(invxor_io_in_key_0_2),
    .io_in_key_0_3(invxor_io_in_key_0_3),
    .io_in_key_1_0(invxor_io_in_key_1_0),
    .io_in_key_1_1(invxor_io_in_key_1_1),
    .io_in_key_1_2(invxor_io_in_key_1_2),
    .io_in_key_1_3(invxor_io_in_key_1_3),
    .io_in_key_2_0(invxor_io_in_key_2_0),
    .io_in_key_2_1(invxor_io_in_key_2_1),
    .io_in_key_2_2(invxor_io_in_key_2_2),
    .io_in_key_2_3(invxor_io_in_key_2_3),
    .io_in_key_3_0(invxor_io_in_key_3_0),
    .io_in_key_3_1(invxor_io_in_key_3_1),
    .io_in_key_3_2(invxor_io_in_key_3_2),
    .io_in_key_3_3(invxor_io_in_key_3_3)
  );
  AES_InvMixColumns invmix ( // @[AES_PipelinedElasticBuffer.scala 189:22]
    .io_out_state_0_0(invmix_io_out_state_0_0),
    .io_out_state_0_1(invmix_io_out_state_0_1),
    .io_out_state_0_2(invmix_io_out_state_0_2),
    .io_out_state_0_3(invmix_io_out_state_0_3),
    .io_out_state_1_0(invmix_io_out_state_1_0),
    .io_out_state_1_1(invmix_io_out_state_1_1),
    .io_out_state_1_2(invmix_io_out_state_1_2),
    .io_out_state_1_3(invmix_io_out_state_1_3),
    .io_out_state_2_0(invmix_io_out_state_2_0),
    .io_out_state_2_1(invmix_io_out_state_2_1),
    .io_out_state_2_2(invmix_io_out_state_2_2),
    .io_out_state_2_3(invmix_io_out_state_2_3),
    .io_out_state_3_0(invmix_io_out_state_3_0),
    .io_out_state_3_1(invmix_io_out_state_3_1),
    .io_out_state_3_2(invmix_io_out_state_3_2),
    .io_out_state_3_3(invmix_io_out_state_3_3),
    .io_in_state_0_0(invmix_io_in_state_0_0),
    .io_in_state_0_1(invmix_io_in_state_0_1),
    .io_in_state_0_2(invmix_io_in_state_0_2),
    .io_in_state_0_3(invmix_io_in_state_0_3),
    .io_in_state_1_0(invmix_io_in_state_1_0),
    .io_in_state_1_1(invmix_io_in_state_1_1),
    .io_in_state_1_2(invmix_io_in_state_1_2),
    .io_in_state_1_3(invmix_io_in_state_1_3),
    .io_in_state_2_0(invmix_io_in_state_2_0),
    .io_in_state_2_1(invmix_io_in_state_2_1),
    .io_in_state_2_2(invmix_io_in_state_2_2),
    .io_in_state_2_3(invmix_io_in_state_2_3),
    .io_in_state_3_0(invmix_io_in_state_3_0),
    .io_in_state_3_1(invmix_io_in_state_3_1),
    .io_in_state_3_2(invmix_io_in_state_3_2),
    .io_in_state_3_3(invmix_io_in_state_3_3)
  );
  AES_InvShiftRows invshift ( // @[AES_PipelinedElasticBuffer.scala 192:24]
    .io_out_state_0_0(invshift_io_out_state_0_0),
    .io_out_state_0_1(invshift_io_out_state_0_1),
    .io_out_state_0_2(invshift_io_out_state_0_2),
    .io_out_state_0_3(invshift_io_out_state_0_3),
    .io_out_state_1_0(invshift_io_out_state_1_0),
    .io_out_state_1_1(invshift_io_out_state_1_1),
    .io_out_state_1_2(invshift_io_out_state_1_2),
    .io_out_state_1_3(invshift_io_out_state_1_3),
    .io_out_state_2_0(invshift_io_out_state_2_0),
    .io_out_state_2_1(invshift_io_out_state_2_1),
    .io_out_state_2_2(invshift_io_out_state_2_2),
    .io_out_state_2_3(invshift_io_out_state_2_3),
    .io_out_state_3_0(invshift_io_out_state_3_0),
    .io_out_state_3_1(invshift_io_out_state_3_1),
    .io_out_state_3_2(invshift_io_out_state_3_2),
    .io_out_state_3_3(invshift_io_out_state_3_3),
    .io_in_state_0_0(invshift_io_in_state_0_0),
    .io_in_state_0_1(invshift_io_in_state_0_1),
    .io_in_state_0_2(invshift_io_in_state_0_2),
    .io_in_state_0_3(invshift_io_in_state_0_3),
    .io_in_state_1_0(invshift_io_in_state_1_0),
    .io_in_state_1_1(invshift_io_in_state_1_1),
    .io_in_state_1_2(invshift_io_in_state_1_2),
    .io_in_state_1_3(invshift_io_in_state_1_3),
    .io_in_state_2_0(invshift_io_in_state_2_0),
    .io_in_state_2_1(invshift_io_in_state_2_1),
    .io_in_state_2_2(invshift_io_in_state_2_2),
    .io_in_state_2_3(invshift_io_in_state_2_3),
    .io_in_state_3_0(invshift_io_in_state_3_0),
    .io_in_state_3_1(invshift_io_in_state_3_1),
    .io_in_state_3_2(invshift_io_in_state_3_2),
    .io_in_state_3_3(invshift_io_in_state_3_3)
  );
  AES_InvSubBytes invsub ( // @[AES_PipelinedElasticBuffer.scala 199:22]
    .io_out_state_0_0(invsub_io_out_state_0_0),
    .io_out_state_0_1(invsub_io_out_state_0_1),
    .io_out_state_0_2(invsub_io_out_state_0_2),
    .io_out_state_0_3(invsub_io_out_state_0_3),
    .io_out_state_1_0(invsub_io_out_state_1_0),
    .io_out_state_1_1(invsub_io_out_state_1_1),
    .io_out_state_1_2(invsub_io_out_state_1_2),
    .io_out_state_1_3(invsub_io_out_state_1_3),
    .io_out_state_2_0(invsub_io_out_state_2_0),
    .io_out_state_2_1(invsub_io_out_state_2_1),
    .io_out_state_2_2(invsub_io_out_state_2_2),
    .io_out_state_2_3(invsub_io_out_state_2_3),
    .io_out_state_3_0(invsub_io_out_state_3_0),
    .io_out_state_3_1(invsub_io_out_state_3_1),
    .io_out_state_3_2(invsub_io_out_state_3_2),
    .io_out_state_3_3(invsub_io_out_state_3_3),
    .io_in_state_0_0(invsub_io_in_state_0_0),
    .io_in_state_0_1(invsub_io_in_state_0_1),
    .io_in_state_0_2(invsub_io_in_state_0_2),
    .io_in_state_0_3(invsub_io_in_state_0_3),
    .io_in_state_1_0(invsub_io_in_state_1_0),
    .io_in_state_1_1(invsub_io_in_state_1_1),
    .io_in_state_1_2(invsub_io_in_state_1_2),
    .io_in_state_1_3(invsub_io_in_state_1_3),
    .io_in_state_2_0(invsub_io_in_state_2_0),
    .io_in_state_2_1(invsub_io_in_state_2_1),
    .io_in_state_2_2(invsub_io_in_state_2_2),
    .io_in_state_2_3(invsub_io_in_state_2_3),
    .io_in_state_3_0(invsub_io_in_state_3_0),
    .io_in_state_3_1(invsub_io_in_state_3_1),
    .io_in_state_3_2(invsub_io_in_state_3_2),
    .io_in_state_3_3(invsub_io_in_state_3_3)
  );
  AES_GetNewKey_2 key ( // @[AES_PipelinedElasticBuffer.scala 202:19]
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  AES_InvGetNewKey_2 invkey ( // @[AES_PipelinedElasticBuffer.scala 206:22]
    .io_out_key_0_0(invkey_io_out_key_0_0),
    .io_out_key_0_1(invkey_io_out_key_0_1),
    .io_out_key_0_2(invkey_io_out_key_0_2),
    .io_out_key_0_3(invkey_io_out_key_0_3),
    .io_out_key_1_0(invkey_io_out_key_1_0),
    .io_out_key_1_1(invkey_io_out_key_1_1),
    .io_out_key_1_2(invkey_io_out_key_1_2),
    .io_out_key_1_3(invkey_io_out_key_1_3),
    .io_out_key_2_0(invkey_io_out_key_2_0),
    .io_out_key_2_1(invkey_io_out_key_2_1),
    .io_out_key_2_2(invkey_io_out_key_2_2),
    .io_out_key_2_3(invkey_io_out_key_2_3),
    .io_out_key_3_0(invkey_io_out_key_3_0),
    .io_out_key_3_1(invkey_io_out_key_3_1),
    .io_out_key_3_2(invkey_io_out_key_3_2),
    .io_out_key_3_3(invkey_io_out_key_3_3),
    .io_in_key_0_0(invkey_io_in_key_0_0),
    .io_in_key_0_1(invkey_io_in_key_0_1),
    .io_in_key_0_2(invkey_io_in_key_0_2),
    .io_in_key_0_3(invkey_io_in_key_0_3),
    .io_in_key_1_0(invkey_io_in_key_1_0),
    .io_in_key_1_1(invkey_io_in_key_1_1),
    .io_in_key_1_2(invkey_io_in_key_1_2),
    .io_in_key_1_3(invkey_io_in_key_1_3),
    .io_in_key_2_0(invkey_io_in_key_2_0),
    .io_in_key_2_1(invkey_io_in_key_2_1),
    .io_in_key_2_2(invkey_io_in_key_2_2),
    .io_in_key_2_3(invkey_io_in_key_2_3),
    .io_in_key_3_0(invkey_io_in_key_3_0),
    .io_in_key_3_1(invkey_io_in_key_3_1),
    .io_in_key_3_2(invkey_io_in_key_3_2),
    .io_in_key_3_3(invkey_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 151:27]
  assign io_out_bits_state_0_0 = invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_1 = invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_2 = invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_3 = invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_0 = invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_1 = invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_2 = invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_3 = invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_0 = invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_1 = invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_2 = invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_3 = invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_0 = invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_1 = invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_2 = invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_3 = invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_0 = invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_1 = invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_2 = invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_3 = invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_0 = invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_1 = invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_2 = invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_3 = invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_0 = invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_1 = invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_2 = invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_3 = invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_0 = invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_1 = invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_2 = invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_3 = invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 150:18]
  assign xor__io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign sub_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign invxor_io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invmix_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invshift_io_in_state_0_0 = invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_1 = invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_2 = invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_3 = invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_0 = invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_1 = invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_2 = invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_3 = invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_0 = invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_1 = invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_2 = invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_3 = invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_0 = invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_1 = invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_2 = invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_3 = invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invsub_io_in_state_0_0 = invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_1 = invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_2 = invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_3 = invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_0 = invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_1 = invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_2 = invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_3 = invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_0 = invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_1 = invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_2 = invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_3 = invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_0 = invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_1 = invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_2 = invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_3 = invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 146:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 146:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 165:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 159:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_3(
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 237:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 240:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 241:13]
endmodule
module AES_InvGetNewKey_3(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] w4 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w5 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w6 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [31:0] w7 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] w3 = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  wire [31:0] w2 = w6 ^ w5; // @[AES_PipelinedElasticBuffer.scala 301:12]
  wire [31:0] w1 = w5 ^ w4; // @[AES_PipelinedElasticBuffer.scala 302:12]
  wire [31:0] temp = 32'h40000000 ^ sub_io_out; // @[AES_PipelinedElasticBuffer.scala 310:16]
  wire [31:0] w0 = w4 ^ temp; // @[AES_PipelinedElasticBuffer.scala 303:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 305:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 308:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w0[31:24]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_1 = w0[23:16]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_2 = w0[15:8]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_3 = w0[7:0]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_1_0 = w1[31:24]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_1 = w1[23:16]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_2 = w1[15:8]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_3 = w1[7:0]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_2_0 = w2[31:24]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_1 = w2[23:16]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_2 = w2[15:8]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_3 = w2[7:0]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_3_0 = w3[31:24]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_1 = w3[23:16]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_2 = w3[15:8]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_3 = w3[7:0]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign rot_io_in = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 309:13]
endmodule
module AES_ProcessingElement_3(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 146:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:23 AES_PipelinedElasticBuffer.scala 156:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 163:21 AES_PipelinedElasticBuffer.scala 163:21]
  AES_XOR xor_ ( // @[AES_PipelinedElasticBuffer.scala 169:19]
    .io_out_state_0_0(xor__io_out_state_0_0),
    .io_out_state_0_1(xor__io_out_state_0_1),
    .io_out_state_0_2(xor__io_out_state_0_2),
    .io_out_state_0_3(xor__io_out_state_0_3),
    .io_out_state_1_0(xor__io_out_state_1_0),
    .io_out_state_1_1(xor__io_out_state_1_1),
    .io_out_state_1_2(xor__io_out_state_1_2),
    .io_out_state_1_3(xor__io_out_state_1_3),
    .io_out_state_2_0(xor__io_out_state_2_0),
    .io_out_state_2_1(xor__io_out_state_2_1),
    .io_out_state_2_2(xor__io_out_state_2_2),
    .io_out_state_2_3(xor__io_out_state_2_3),
    .io_out_state_3_0(xor__io_out_state_3_0),
    .io_out_state_3_1(xor__io_out_state_3_1),
    .io_out_state_3_2(xor__io_out_state_3_2),
    .io_out_state_3_3(xor__io_out_state_3_3),
    .io_in_state_0_0(xor__io_in_state_0_0),
    .io_in_state_0_1(xor__io_in_state_0_1),
    .io_in_state_0_2(xor__io_in_state_0_2),
    .io_in_state_0_3(xor__io_in_state_0_3),
    .io_in_state_1_0(xor__io_in_state_1_0),
    .io_in_state_1_1(xor__io_in_state_1_1),
    .io_in_state_1_2(xor__io_in_state_1_2),
    .io_in_state_1_3(xor__io_in_state_1_3),
    .io_in_state_2_0(xor__io_in_state_2_0),
    .io_in_state_2_1(xor__io_in_state_2_1),
    .io_in_state_2_2(xor__io_in_state_2_2),
    .io_in_state_2_3(xor__io_in_state_2_3),
    .io_in_state_3_0(xor__io_in_state_3_0),
    .io_in_state_3_1(xor__io_in_state_3_1),
    .io_in_state_3_2(xor__io_in_state_3_2),
    .io_in_state_3_3(xor__io_in_state_3_3),
    .io_in_key_0_0(xor__io_in_key_0_0),
    .io_in_key_0_1(xor__io_in_key_0_1),
    .io_in_key_0_2(xor__io_in_key_0_2),
    .io_in_key_0_3(xor__io_in_key_0_3),
    .io_in_key_1_0(xor__io_in_key_1_0),
    .io_in_key_1_1(xor__io_in_key_1_1),
    .io_in_key_1_2(xor__io_in_key_1_2),
    .io_in_key_1_3(xor__io_in_key_1_3),
    .io_in_key_2_0(xor__io_in_key_2_0),
    .io_in_key_2_1(xor__io_in_key_2_1),
    .io_in_key_2_2(xor__io_in_key_2_2),
    .io_in_key_2_3(xor__io_in_key_2_3),
    .io_in_key_3_0(xor__io_in_key_3_0),
    .io_in_key_3_1(xor__io_in_key_3_1),
    .io_in_key_3_2(xor__io_in_key_3_2),
    .io_in_key_3_3(xor__io_in_key_3_3)
  );
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 174:19]
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_XOR invxor ( // @[AES_PipelinedElasticBuffer.scala 184:22]
    .io_out_state_0_0(invxor_io_out_state_0_0),
    .io_out_state_0_1(invxor_io_out_state_0_1),
    .io_out_state_0_2(invxor_io_out_state_0_2),
    .io_out_state_0_3(invxor_io_out_state_0_3),
    .io_out_state_1_0(invxor_io_out_state_1_0),
    .io_out_state_1_1(invxor_io_out_state_1_1),
    .io_out_state_1_2(invxor_io_out_state_1_2),
    .io_out_state_1_3(invxor_io_out_state_1_3),
    .io_out_state_2_0(invxor_io_out_state_2_0),
    .io_out_state_2_1(invxor_io_out_state_2_1),
    .io_out_state_2_2(invxor_io_out_state_2_2),
    .io_out_state_2_3(invxor_io_out_state_2_3),
    .io_out_state_3_0(invxor_io_out_state_3_0),
    .io_out_state_3_1(invxor_io_out_state_3_1),
    .io_out_state_3_2(invxor_io_out_state_3_2),
    .io_out_state_3_3(invxor_io_out_state_3_3),
    .io_in_state_0_0(invxor_io_in_state_0_0),
    .io_in_state_0_1(invxor_io_in_state_0_1),
    .io_in_state_0_2(invxor_io_in_state_0_2),
    .io_in_state_0_3(invxor_io_in_state_0_3),
    .io_in_state_1_0(invxor_io_in_state_1_0),
    .io_in_state_1_1(invxor_io_in_state_1_1),
    .io_in_state_1_2(invxor_io_in_state_1_2),
    .io_in_state_1_3(invxor_io_in_state_1_3),
    .io_in_state_2_0(invxor_io_in_state_2_0),
    .io_in_state_2_1(invxor_io_in_state_2_1),
    .io_in_state_2_2(invxor_io_in_state_2_2),
    .io_in_state_2_3(invxor_io_in_state_2_3),
    .io_in_state_3_0(invxor_io_in_state_3_0),
    .io_in_state_3_1(invxor_io_in_state_3_1),
    .io_in_state_3_2(invxor_io_in_state_3_2),
    .io_in_state_3_3(invxor_io_in_state_3_3),
    .io_in_key_0_0(invxor_io_in_key_0_0),
    .io_in_key_0_1(invxor_io_in_key_0_1),
    .io_in_key_0_2(invxor_io_in_key_0_2),
    .io_in_key_0_3(invxor_io_in_key_0_3),
    .io_in_key_1_0(invxor_io_in_key_1_0),
    .io_in_key_1_1(invxor_io_in_key_1_1),
    .io_in_key_1_2(invxor_io_in_key_1_2),
    .io_in_key_1_3(invxor_io_in_key_1_3),
    .io_in_key_2_0(invxor_io_in_key_2_0),
    .io_in_key_2_1(invxor_io_in_key_2_1),
    .io_in_key_2_2(invxor_io_in_key_2_2),
    .io_in_key_2_3(invxor_io_in_key_2_3),
    .io_in_key_3_0(invxor_io_in_key_3_0),
    .io_in_key_3_1(invxor_io_in_key_3_1),
    .io_in_key_3_2(invxor_io_in_key_3_2),
    .io_in_key_3_3(invxor_io_in_key_3_3)
  );
  AES_InvMixColumns invmix ( // @[AES_PipelinedElasticBuffer.scala 189:22]
    .io_out_state_0_0(invmix_io_out_state_0_0),
    .io_out_state_0_1(invmix_io_out_state_0_1),
    .io_out_state_0_2(invmix_io_out_state_0_2),
    .io_out_state_0_3(invmix_io_out_state_0_3),
    .io_out_state_1_0(invmix_io_out_state_1_0),
    .io_out_state_1_1(invmix_io_out_state_1_1),
    .io_out_state_1_2(invmix_io_out_state_1_2),
    .io_out_state_1_3(invmix_io_out_state_1_3),
    .io_out_state_2_0(invmix_io_out_state_2_0),
    .io_out_state_2_1(invmix_io_out_state_2_1),
    .io_out_state_2_2(invmix_io_out_state_2_2),
    .io_out_state_2_3(invmix_io_out_state_2_3),
    .io_out_state_3_0(invmix_io_out_state_3_0),
    .io_out_state_3_1(invmix_io_out_state_3_1),
    .io_out_state_3_2(invmix_io_out_state_3_2),
    .io_out_state_3_3(invmix_io_out_state_3_3),
    .io_in_state_0_0(invmix_io_in_state_0_0),
    .io_in_state_0_1(invmix_io_in_state_0_1),
    .io_in_state_0_2(invmix_io_in_state_0_2),
    .io_in_state_0_3(invmix_io_in_state_0_3),
    .io_in_state_1_0(invmix_io_in_state_1_0),
    .io_in_state_1_1(invmix_io_in_state_1_1),
    .io_in_state_1_2(invmix_io_in_state_1_2),
    .io_in_state_1_3(invmix_io_in_state_1_3),
    .io_in_state_2_0(invmix_io_in_state_2_0),
    .io_in_state_2_1(invmix_io_in_state_2_1),
    .io_in_state_2_2(invmix_io_in_state_2_2),
    .io_in_state_2_3(invmix_io_in_state_2_3),
    .io_in_state_3_0(invmix_io_in_state_3_0),
    .io_in_state_3_1(invmix_io_in_state_3_1),
    .io_in_state_3_2(invmix_io_in_state_3_2),
    .io_in_state_3_3(invmix_io_in_state_3_3)
  );
  AES_InvShiftRows invshift ( // @[AES_PipelinedElasticBuffer.scala 192:24]
    .io_out_state_0_0(invshift_io_out_state_0_0),
    .io_out_state_0_1(invshift_io_out_state_0_1),
    .io_out_state_0_2(invshift_io_out_state_0_2),
    .io_out_state_0_3(invshift_io_out_state_0_3),
    .io_out_state_1_0(invshift_io_out_state_1_0),
    .io_out_state_1_1(invshift_io_out_state_1_1),
    .io_out_state_1_2(invshift_io_out_state_1_2),
    .io_out_state_1_3(invshift_io_out_state_1_3),
    .io_out_state_2_0(invshift_io_out_state_2_0),
    .io_out_state_2_1(invshift_io_out_state_2_1),
    .io_out_state_2_2(invshift_io_out_state_2_2),
    .io_out_state_2_3(invshift_io_out_state_2_3),
    .io_out_state_3_0(invshift_io_out_state_3_0),
    .io_out_state_3_1(invshift_io_out_state_3_1),
    .io_out_state_3_2(invshift_io_out_state_3_2),
    .io_out_state_3_3(invshift_io_out_state_3_3),
    .io_in_state_0_0(invshift_io_in_state_0_0),
    .io_in_state_0_1(invshift_io_in_state_0_1),
    .io_in_state_0_2(invshift_io_in_state_0_2),
    .io_in_state_0_3(invshift_io_in_state_0_3),
    .io_in_state_1_0(invshift_io_in_state_1_0),
    .io_in_state_1_1(invshift_io_in_state_1_1),
    .io_in_state_1_2(invshift_io_in_state_1_2),
    .io_in_state_1_3(invshift_io_in_state_1_3),
    .io_in_state_2_0(invshift_io_in_state_2_0),
    .io_in_state_2_1(invshift_io_in_state_2_1),
    .io_in_state_2_2(invshift_io_in_state_2_2),
    .io_in_state_2_3(invshift_io_in_state_2_3),
    .io_in_state_3_0(invshift_io_in_state_3_0),
    .io_in_state_3_1(invshift_io_in_state_3_1),
    .io_in_state_3_2(invshift_io_in_state_3_2),
    .io_in_state_3_3(invshift_io_in_state_3_3)
  );
  AES_InvSubBytes invsub ( // @[AES_PipelinedElasticBuffer.scala 199:22]
    .io_out_state_0_0(invsub_io_out_state_0_0),
    .io_out_state_0_1(invsub_io_out_state_0_1),
    .io_out_state_0_2(invsub_io_out_state_0_2),
    .io_out_state_0_3(invsub_io_out_state_0_3),
    .io_out_state_1_0(invsub_io_out_state_1_0),
    .io_out_state_1_1(invsub_io_out_state_1_1),
    .io_out_state_1_2(invsub_io_out_state_1_2),
    .io_out_state_1_3(invsub_io_out_state_1_3),
    .io_out_state_2_0(invsub_io_out_state_2_0),
    .io_out_state_2_1(invsub_io_out_state_2_1),
    .io_out_state_2_2(invsub_io_out_state_2_2),
    .io_out_state_2_3(invsub_io_out_state_2_3),
    .io_out_state_3_0(invsub_io_out_state_3_0),
    .io_out_state_3_1(invsub_io_out_state_3_1),
    .io_out_state_3_2(invsub_io_out_state_3_2),
    .io_out_state_3_3(invsub_io_out_state_3_3),
    .io_in_state_0_0(invsub_io_in_state_0_0),
    .io_in_state_0_1(invsub_io_in_state_0_1),
    .io_in_state_0_2(invsub_io_in_state_0_2),
    .io_in_state_0_3(invsub_io_in_state_0_3),
    .io_in_state_1_0(invsub_io_in_state_1_0),
    .io_in_state_1_1(invsub_io_in_state_1_1),
    .io_in_state_1_2(invsub_io_in_state_1_2),
    .io_in_state_1_3(invsub_io_in_state_1_3),
    .io_in_state_2_0(invsub_io_in_state_2_0),
    .io_in_state_2_1(invsub_io_in_state_2_1),
    .io_in_state_2_2(invsub_io_in_state_2_2),
    .io_in_state_2_3(invsub_io_in_state_2_3),
    .io_in_state_3_0(invsub_io_in_state_3_0),
    .io_in_state_3_1(invsub_io_in_state_3_1),
    .io_in_state_3_2(invsub_io_in_state_3_2),
    .io_in_state_3_3(invsub_io_in_state_3_3)
  );
  AES_GetNewKey_3 key ( // @[AES_PipelinedElasticBuffer.scala 202:19]
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  AES_InvGetNewKey_3 invkey ( // @[AES_PipelinedElasticBuffer.scala 206:22]
    .io_out_key_0_0(invkey_io_out_key_0_0),
    .io_out_key_0_1(invkey_io_out_key_0_1),
    .io_out_key_0_2(invkey_io_out_key_0_2),
    .io_out_key_0_3(invkey_io_out_key_0_3),
    .io_out_key_1_0(invkey_io_out_key_1_0),
    .io_out_key_1_1(invkey_io_out_key_1_1),
    .io_out_key_1_2(invkey_io_out_key_1_2),
    .io_out_key_1_3(invkey_io_out_key_1_3),
    .io_out_key_2_0(invkey_io_out_key_2_0),
    .io_out_key_2_1(invkey_io_out_key_2_1),
    .io_out_key_2_2(invkey_io_out_key_2_2),
    .io_out_key_2_3(invkey_io_out_key_2_3),
    .io_out_key_3_0(invkey_io_out_key_3_0),
    .io_out_key_3_1(invkey_io_out_key_3_1),
    .io_out_key_3_2(invkey_io_out_key_3_2),
    .io_out_key_3_3(invkey_io_out_key_3_3),
    .io_in_key_0_0(invkey_io_in_key_0_0),
    .io_in_key_0_1(invkey_io_in_key_0_1),
    .io_in_key_0_2(invkey_io_in_key_0_2),
    .io_in_key_0_3(invkey_io_in_key_0_3),
    .io_in_key_1_0(invkey_io_in_key_1_0),
    .io_in_key_1_1(invkey_io_in_key_1_1),
    .io_in_key_1_2(invkey_io_in_key_1_2),
    .io_in_key_1_3(invkey_io_in_key_1_3),
    .io_in_key_2_0(invkey_io_in_key_2_0),
    .io_in_key_2_1(invkey_io_in_key_2_1),
    .io_in_key_2_2(invkey_io_in_key_2_2),
    .io_in_key_2_3(invkey_io_in_key_2_3),
    .io_in_key_3_0(invkey_io_in_key_3_0),
    .io_in_key_3_1(invkey_io_in_key_3_1),
    .io_in_key_3_2(invkey_io_in_key_3_2),
    .io_in_key_3_3(invkey_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 151:27]
  assign io_out_bits_state_0_0 = invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_1 = invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_2 = invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_3 = invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_0 = invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_1 = invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_2 = invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_3 = invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_0 = invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_1 = invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_2 = invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_3 = invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_0 = invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_1 = invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_2 = invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_3 = invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_0 = invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_1 = invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_2 = invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_3 = invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_0 = invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_1 = invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_2 = invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_3 = invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_0 = invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_1 = invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_2 = invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_3 = invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_0 = invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_1 = invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_2 = invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_3 = invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 150:18]
  assign xor__io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign sub_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign invxor_io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invmix_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invshift_io_in_state_0_0 = invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_1 = invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_2 = invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_3 = invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_0 = invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_1 = invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_2 = invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_3 = invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_0 = invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_1 = invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_2 = invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_3 = invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_0 = invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_1 = invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_2 = invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_3 = invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invsub_io_in_state_0_0 = invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_1 = invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_2 = invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_3 = invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_0 = invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_1 = invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_2 = invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_3 = invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_0 = invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_1 = invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_2 = invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_3 = invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_0 = invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_1 = invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_2 = invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_3 = invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 146:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 146:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 165:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 159:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_4(
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 237:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 240:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 241:13]
endmodule
module AES_InvGetNewKey_4(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] w4 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w5 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w6 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [31:0] w7 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] w3 = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  wire [31:0] w2 = w6 ^ w5; // @[AES_PipelinedElasticBuffer.scala 301:12]
  wire [31:0] w1 = w5 ^ w4; // @[AES_PipelinedElasticBuffer.scala 302:12]
  wire [31:0] temp = 32'h20000000 ^ sub_io_out; // @[AES_PipelinedElasticBuffer.scala 310:16]
  wire [31:0] w0 = w4 ^ temp; // @[AES_PipelinedElasticBuffer.scala 303:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 305:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 308:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w0[31:24]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_1 = w0[23:16]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_2 = w0[15:8]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_3 = w0[7:0]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_1_0 = w1[31:24]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_1 = w1[23:16]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_2 = w1[15:8]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_3 = w1[7:0]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_2_0 = w2[31:24]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_1 = w2[23:16]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_2 = w2[15:8]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_3 = w2[7:0]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_3_0 = w3[31:24]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_1 = w3[23:16]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_2 = w3[15:8]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_3 = w3[7:0]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign rot_io_in = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 309:13]
endmodule
module AES_ProcessingElement_4(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 146:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:23 AES_PipelinedElasticBuffer.scala 156:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 163:21 AES_PipelinedElasticBuffer.scala 163:21]
  AES_XOR xor_ ( // @[AES_PipelinedElasticBuffer.scala 169:19]
    .io_out_state_0_0(xor__io_out_state_0_0),
    .io_out_state_0_1(xor__io_out_state_0_1),
    .io_out_state_0_2(xor__io_out_state_0_2),
    .io_out_state_0_3(xor__io_out_state_0_3),
    .io_out_state_1_0(xor__io_out_state_1_0),
    .io_out_state_1_1(xor__io_out_state_1_1),
    .io_out_state_1_2(xor__io_out_state_1_2),
    .io_out_state_1_3(xor__io_out_state_1_3),
    .io_out_state_2_0(xor__io_out_state_2_0),
    .io_out_state_2_1(xor__io_out_state_2_1),
    .io_out_state_2_2(xor__io_out_state_2_2),
    .io_out_state_2_3(xor__io_out_state_2_3),
    .io_out_state_3_0(xor__io_out_state_3_0),
    .io_out_state_3_1(xor__io_out_state_3_1),
    .io_out_state_3_2(xor__io_out_state_3_2),
    .io_out_state_3_3(xor__io_out_state_3_3),
    .io_in_state_0_0(xor__io_in_state_0_0),
    .io_in_state_0_1(xor__io_in_state_0_1),
    .io_in_state_0_2(xor__io_in_state_0_2),
    .io_in_state_0_3(xor__io_in_state_0_3),
    .io_in_state_1_0(xor__io_in_state_1_0),
    .io_in_state_1_1(xor__io_in_state_1_1),
    .io_in_state_1_2(xor__io_in_state_1_2),
    .io_in_state_1_3(xor__io_in_state_1_3),
    .io_in_state_2_0(xor__io_in_state_2_0),
    .io_in_state_2_1(xor__io_in_state_2_1),
    .io_in_state_2_2(xor__io_in_state_2_2),
    .io_in_state_2_3(xor__io_in_state_2_3),
    .io_in_state_3_0(xor__io_in_state_3_0),
    .io_in_state_3_1(xor__io_in_state_3_1),
    .io_in_state_3_2(xor__io_in_state_3_2),
    .io_in_state_3_3(xor__io_in_state_3_3),
    .io_in_key_0_0(xor__io_in_key_0_0),
    .io_in_key_0_1(xor__io_in_key_0_1),
    .io_in_key_0_2(xor__io_in_key_0_2),
    .io_in_key_0_3(xor__io_in_key_0_3),
    .io_in_key_1_0(xor__io_in_key_1_0),
    .io_in_key_1_1(xor__io_in_key_1_1),
    .io_in_key_1_2(xor__io_in_key_1_2),
    .io_in_key_1_3(xor__io_in_key_1_3),
    .io_in_key_2_0(xor__io_in_key_2_0),
    .io_in_key_2_1(xor__io_in_key_2_1),
    .io_in_key_2_2(xor__io_in_key_2_2),
    .io_in_key_2_3(xor__io_in_key_2_3),
    .io_in_key_3_0(xor__io_in_key_3_0),
    .io_in_key_3_1(xor__io_in_key_3_1),
    .io_in_key_3_2(xor__io_in_key_3_2),
    .io_in_key_3_3(xor__io_in_key_3_3)
  );
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 174:19]
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_XOR invxor ( // @[AES_PipelinedElasticBuffer.scala 184:22]
    .io_out_state_0_0(invxor_io_out_state_0_0),
    .io_out_state_0_1(invxor_io_out_state_0_1),
    .io_out_state_0_2(invxor_io_out_state_0_2),
    .io_out_state_0_3(invxor_io_out_state_0_3),
    .io_out_state_1_0(invxor_io_out_state_1_0),
    .io_out_state_1_1(invxor_io_out_state_1_1),
    .io_out_state_1_2(invxor_io_out_state_1_2),
    .io_out_state_1_3(invxor_io_out_state_1_3),
    .io_out_state_2_0(invxor_io_out_state_2_0),
    .io_out_state_2_1(invxor_io_out_state_2_1),
    .io_out_state_2_2(invxor_io_out_state_2_2),
    .io_out_state_2_3(invxor_io_out_state_2_3),
    .io_out_state_3_0(invxor_io_out_state_3_0),
    .io_out_state_3_1(invxor_io_out_state_3_1),
    .io_out_state_3_2(invxor_io_out_state_3_2),
    .io_out_state_3_3(invxor_io_out_state_3_3),
    .io_in_state_0_0(invxor_io_in_state_0_0),
    .io_in_state_0_1(invxor_io_in_state_0_1),
    .io_in_state_0_2(invxor_io_in_state_0_2),
    .io_in_state_0_3(invxor_io_in_state_0_3),
    .io_in_state_1_0(invxor_io_in_state_1_0),
    .io_in_state_1_1(invxor_io_in_state_1_1),
    .io_in_state_1_2(invxor_io_in_state_1_2),
    .io_in_state_1_3(invxor_io_in_state_1_3),
    .io_in_state_2_0(invxor_io_in_state_2_0),
    .io_in_state_2_1(invxor_io_in_state_2_1),
    .io_in_state_2_2(invxor_io_in_state_2_2),
    .io_in_state_2_3(invxor_io_in_state_2_3),
    .io_in_state_3_0(invxor_io_in_state_3_0),
    .io_in_state_3_1(invxor_io_in_state_3_1),
    .io_in_state_3_2(invxor_io_in_state_3_2),
    .io_in_state_3_3(invxor_io_in_state_3_3),
    .io_in_key_0_0(invxor_io_in_key_0_0),
    .io_in_key_0_1(invxor_io_in_key_0_1),
    .io_in_key_0_2(invxor_io_in_key_0_2),
    .io_in_key_0_3(invxor_io_in_key_0_3),
    .io_in_key_1_0(invxor_io_in_key_1_0),
    .io_in_key_1_1(invxor_io_in_key_1_1),
    .io_in_key_1_2(invxor_io_in_key_1_2),
    .io_in_key_1_3(invxor_io_in_key_1_3),
    .io_in_key_2_0(invxor_io_in_key_2_0),
    .io_in_key_2_1(invxor_io_in_key_2_1),
    .io_in_key_2_2(invxor_io_in_key_2_2),
    .io_in_key_2_3(invxor_io_in_key_2_3),
    .io_in_key_3_0(invxor_io_in_key_3_0),
    .io_in_key_3_1(invxor_io_in_key_3_1),
    .io_in_key_3_2(invxor_io_in_key_3_2),
    .io_in_key_3_3(invxor_io_in_key_3_3)
  );
  AES_InvMixColumns invmix ( // @[AES_PipelinedElasticBuffer.scala 189:22]
    .io_out_state_0_0(invmix_io_out_state_0_0),
    .io_out_state_0_1(invmix_io_out_state_0_1),
    .io_out_state_0_2(invmix_io_out_state_0_2),
    .io_out_state_0_3(invmix_io_out_state_0_3),
    .io_out_state_1_0(invmix_io_out_state_1_0),
    .io_out_state_1_1(invmix_io_out_state_1_1),
    .io_out_state_1_2(invmix_io_out_state_1_2),
    .io_out_state_1_3(invmix_io_out_state_1_3),
    .io_out_state_2_0(invmix_io_out_state_2_0),
    .io_out_state_2_1(invmix_io_out_state_2_1),
    .io_out_state_2_2(invmix_io_out_state_2_2),
    .io_out_state_2_3(invmix_io_out_state_2_3),
    .io_out_state_3_0(invmix_io_out_state_3_0),
    .io_out_state_3_1(invmix_io_out_state_3_1),
    .io_out_state_3_2(invmix_io_out_state_3_2),
    .io_out_state_3_3(invmix_io_out_state_3_3),
    .io_in_state_0_0(invmix_io_in_state_0_0),
    .io_in_state_0_1(invmix_io_in_state_0_1),
    .io_in_state_0_2(invmix_io_in_state_0_2),
    .io_in_state_0_3(invmix_io_in_state_0_3),
    .io_in_state_1_0(invmix_io_in_state_1_0),
    .io_in_state_1_1(invmix_io_in_state_1_1),
    .io_in_state_1_2(invmix_io_in_state_1_2),
    .io_in_state_1_3(invmix_io_in_state_1_3),
    .io_in_state_2_0(invmix_io_in_state_2_0),
    .io_in_state_2_1(invmix_io_in_state_2_1),
    .io_in_state_2_2(invmix_io_in_state_2_2),
    .io_in_state_2_3(invmix_io_in_state_2_3),
    .io_in_state_3_0(invmix_io_in_state_3_0),
    .io_in_state_3_1(invmix_io_in_state_3_1),
    .io_in_state_3_2(invmix_io_in_state_3_2),
    .io_in_state_3_3(invmix_io_in_state_3_3)
  );
  AES_InvShiftRows invshift ( // @[AES_PipelinedElasticBuffer.scala 192:24]
    .io_out_state_0_0(invshift_io_out_state_0_0),
    .io_out_state_0_1(invshift_io_out_state_0_1),
    .io_out_state_0_2(invshift_io_out_state_0_2),
    .io_out_state_0_3(invshift_io_out_state_0_3),
    .io_out_state_1_0(invshift_io_out_state_1_0),
    .io_out_state_1_1(invshift_io_out_state_1_1),
    .io_out_state_1_2(invshift_io_out_state_1_2),
    .io_out_state_1_3(invshift_io_out_state_1_3),
    .io_out_state_2_0(invshift_io_out_state_2_0),
    .io_out_state_2_1(invshift_io_out_state_2_1),
    .io_out_state_2_2(invshift_io_out_state_2_2),
    .io_out_state_2_3(invshift_io_out_state_2_3),
    .io_out_state_3_0(invshift_io_out_state_3_0),
    .io_out_state_3_1(invshift_io_out_state_3_1),
    .io_out_state_3_2(invshift_io_out_state_3_2),
    .io_out_state_3_3(invshift_io_out_state_3_3),
    .io_in_state_0_0(invshift_io_in_state_0_0),
    .io_in_state_0_1(invshift_io_in_state_0_1),
    .io_in_state_0_2(invshift_io_in_state_0_2),
    .io_in_state_0_3(invshift_io_in_state_0_3),
    .io_in_state_1_0(invshift_io_in_state_1_0),
    .io_in_state_1_1(invshift_io_in_state_1_1),
    .io_in_state_1_2(invshift_io_in_state_1_2),
    .io_in_state_1_3(invshift_io_in_state_1_3),
    .io_in_state_2_0(invshift_io_in_state_2_0),
    .io_in_state_2_1(invshift_io_in_state_2_1),
    .io_in_state_2_2(invshift_io_in_state_2_2),
    .io_in_state_2_3(invshift_io_in_state_2_3),
    .io_in_state_3_0(invshift_io_in_state_3_0),
    .io_in_state_3_1(invshift_io_in_state_3_1),
    .io_in_state_3_2(invshift_io_in_state_3_2),
    .io_in_state_3_3(invshift_io_in_state_3_3)
  );
  AES_InvSubBytes invsub ( // @[AES_PipelinedElasticBuffer.scala 199:22]
    .io_out_state_0_0(invsub_io_out_state_0_0),
    .io_out_state_0_1(invsub_io_out_state_0_1),
    .io_out_state_0_2(invsub_io_out_state_0_2),
    .io_out_state_0_3(invsub_io_out_state_0_3),
    .io_out_state_1_0(invsub_io_out_state_1_0),
    .io_out_state_1_1(invsub_io_out_state_1_1),
    .io_out_state_1_2(invsub_io_out_state_1_2),
    .io_out_state_1_3(invsub_io_out_state_1_3),
    .io_out_state_2_0(invsub_io_out_state_2_0),
    .io_out_state_2_1(invsub_io_out_state_2_1),
    .io_out_state_2_2(invsub_io_out_state_2_2),
    .io_out_state_2_3(invsub_io_out_state_2_3),
    .io_out_state_3_0(invsub_io_out_state_3_0),
    .io_out_state_3_1(invsub_io_out_state_3_1),
    .io_out_state_3_2(invsub_io_out_state_3_2),
    .io_out_state_3_3(invsub_io_out_state_3_3),
    .io_in_state_0_0(invsub_io_in_state_0_0),
    .io_in_state_0_1(invsub_io_in_state_0_1),
    .io_in_state_0_2(invsub_io_in_state_0_2),
    .io_in_state_0_3(invsub_io_in_state_0_3),
    .io_in_state_1_0(invsub_io_in_state_1_0),
    .io_in_state_1_1(invsub_io_in_state_1_1),
    .io_in_state_1_2(invsub_io_in_state_1_2),
    .io_in_state_1_3(invsub_io_in_state_1_3),
    .io_in_state_2_0(invsub_io_in_state_2_0),
    .io_in_state_2_1(invsub_io_in_state_2_1),
    .io_in_state_2_2(invsub_io_in_state_2_2),
    .io_in_state_2_3(invsub_io_in_state_2_3),
    .io_in_state_3_0(invsub_io_in_state_3_0),
    .io_in_state_3_1(invsub_io_in_state_3_1),
    .io_in_state_3_2(invsub_io_in_state_3_2),
    .io_in_state_3_3(invsub_io_in_state_3_3)
  );
  AES_GetNewKey_4 key ( // @[AES_PipelinedElasticBuffer.scala 202:19]
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  AES_InvGetNewKey_4 invkey ( // @[AES_PipelinedElasticBuffer.scala 206:22]
    .io_out_key_0_0(invkey_io_out_key_0_0),
    .io_out_key_0_1(invkey_io_out_key_0_1),
    .io_out_key_0_2(invkey_io_out_key_0_2),
    .io_out_key_0_3(invkey_io_out_key_0_3),
    .io_out_key_1_0(invkey_io_out_key_1_0),
    .io_out_key_1_1(invkey_io_out_key_1_1),
    .io_out_key_1_2(invkey_io_out_key_1_2),
    .io_out_key_1_3(invkey_io_out_key_1_3),
    .io_out_key_2_0(invkey_io_out_key_2_0),
    .io_out_key_2_1(invkey_io_out_key_2_1),
    .io_out_key_2_2(invkey_io_out_key_2_2),
    .io_out_key_2_3(invkey_io_out_key_2_3),
    .io_out_key_3_0(invkey_io_out_key_3_0),
    .io_out_key_3_1(invkey_io_out_key_3_1),
    .io_out_key_3_2(invkey_io_out_key_3_2),
    .io_out_key_3_3(invkey_io_out_key_3_3),
    .io_in_key_0_0(invkey_io_in_key_0_0),
    .io_in_key_0_1(invkey_io_in_key_0_1),
    .io_in_key_0_2(invkey_io_in_key_0_2),
    .io_in_key_0_3(invkey_io_in_key_0_3),
    .io_in_key_1_0(invkey_io_in_key_1_0),
    .io_in_key_1_1(invkey_io_in_key_1_1),
    .io_in_key_1_2(invkey_io_in_key_1_2),
    .io_in_key_1_3(invkey_io_in_key_1_3),
    .io_in_key_2_0(invkey_io_in_key_2_0),
    .io_in_key_2_1(invkey_io_in_key_2_1),
    .io_in_key_2_2(invkey_io_in_key_2_2),
    .io_in_key_2_3(invkey_io_in_key_2_3),
    .io_in_key_3_0(invkey_io_in_key_3_0),
    .io_in_key_3_1(invkey_io_in_key_3_1),
    .io_in_key_3_2(invkey_io_in_key_3_2),
    .io_in_key_3_3(invkey_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 151:27]
  assign io_out_bits_state_0_0 = invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_1 = invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_2 = invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_3 = invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_0 = invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_1 = invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_2 = invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_3 = invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_0 = invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_1 = invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_2 = invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_3 = invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_0 = invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_1 = invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_2 = invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_3 = invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_0 = invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_1 = invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_2 = invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_3 = invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_0 = invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_1 = invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_2 = invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_3 = invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_0 = invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_1 = invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_2 = invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_3 = invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_0 = invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_1 = invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_2 = invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_3 = invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 150:18]
  assign xor__io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign sub_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign invxor_io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invmix_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invshift_io_in_state_0_0 = invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_1 = invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_2 = invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_3 = invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_0 = invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_1 = invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_2 = invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_3 = invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_0 = invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_1 = invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_2 = invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_3 = invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_0 = invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_1 = invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_2 = invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_3 = invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invsub_io_in_state_0_0 = invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_1 = invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_2 = invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_3 = invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_0 = invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_1 = invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_2 = invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_3 = invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_0 = invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_1 = invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_2 = invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_3 = invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_0 = invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_1 = invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_2 = invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_3 = invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 146:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 146:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 165:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 159:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_5(
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 237:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 240:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 241:13]
endmodule
module AES_InvGetNewKey_5(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] w4 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w5 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w6 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [31:0] w7 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] w3 = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  wire [31:0] w2 = w6 ^ w5; // @[AES_PipelinedElasticBuffer.scala 301:12]
  wire [31:0] w1 = w5 ^ w4; // @[AES_PipelinedElasticBuffer.scala 302:12]
  wire [31:0] temp = 32'h10000000 ^ sub_io_out; // @[AES_PipelinedElasticBuffer.scala 310:16]
  wire [31:0] w0 = w4 ^ temp; // @[AES_PipelinedElasticBuffer.scala 303:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 305:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 308:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w0[31:24]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_1 = w0[23:16]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_2 = w0[15:8]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_3 = w0[7:0]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_1_0 = w1[31:24]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_1 = w1[23:16]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_2 = w1[15:8]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_3 = w1[7:0]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_2_0 = w2[31:24]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_1 = w2[23:16]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_2 = w2[15:8]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_3 = w2[7:0]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_3_0 = w3[31:24]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_1 = w3[23:16]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_2 = w3[15:8]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_3 = w3[7:0]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign rot_io_in = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 309:13]
endmodule
module AES_ProcessingElement_5(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 146:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:23 AES_PipelinedElasticBuffer.scala 156:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 163:21 AES_PipelinedElasticBuffer.scala 163:21]
  AES_XOR xor_ ( // @[AES_PipelinedElasticBuffer.scala 169:19]
    .io_out_state_0_0(xor__io_out_state_0_0),
    .io_out_state_0_1(xor__io_out_state_0_1),
    .io_out_state_0_2(xor__io_out_state_0_2),
    .io_out_state_0_3(xor__io_out_state_0_3),
    .io_out_state_1_0(xor__io_out_state_1_0),
    .io_out_state_1_1(xor__io_out_state_1_1),
    .io_out_state_1_2(xor__io_out_state_1_2),
    .io_out_state_1_3(xor__io_out_state_1_3),
    .io_out_state_2_0(xor__io_out_state_2_0),
    .io_out_state_2_1(xor__io_out_state_2_1),
    .io_out_state_2_2(xor__io_out_state_2_2),
    .io_out_state_2_3(xor__io_out_state_2_3),
    .io_out_state_3_0(xor__io_out_state_3_0),
    .io_out_state_3_1(xor__io_out_state_3_1),
    .io_out_state_3_2(xor__io_out_state_3_2),
    .io_out_state_3_3(xor__io_out_state_3_3),
    .io_in_state_0_0(xor__io_in_state_0_0),
    .io_in_state_0_1(xor__io_in_state_0_1),
    .io_in_state_0_2(xor__io_in_state_0_2),
    .io_in_state_0_3(xor__io_in_state_0_3),
    .io_in_state_1_0(xor__io_in_state_1_0),
    .io_in_state_1_1(xor__io_in_state_1_1),
    .io_in_state_1_2(xor__io_in_state_1_2),
    .io_in_state_1_3(xor__io_in_state_1_3),
    .io_in_state_2_0(xor__io_in_state_2_0),
    .io_in_state_2_1(xor__io_in_state_2_1),
    .io_in_state_2_2(xor__io_in_state_2_2),
    .io_in_state_2_3(xor__io_in_state_2_3),
    .io_in_state_3_0(xor__io_in_state_3_0),
    .io_in_state_3_1(xor__io_in_state_3_1),
    .io_in_state_3_2(xor__io_in_state_3_2),
    .io_in_state_3_3(xor__io_in_state_3_3),
    .io_in_key_0_0(xor__io_in_key_0_0),
    .io_in_key_0_1(xor__io_in_key_0_1),
    .io_in_key_0_2(xor__io_in_key_0_2),
    .io_in_key_0_3(xor__io_in_key_0_3),
    .io_in_key_1_0(xor__io_in_key_1_0),
    .io_in_key_1_1(xor__io_in_key_1_1),
    .io_in_key_1_2(xor__io_in_key_1_2),
    .io_in_key_1_3(xor__io_in_key_1_3),
    .io_in_key_2_0(xor__io_in_key_2_0),
    .io_in_key_2_1(xor__io_in_key_2_1),
    .io_in_key_2_2(xor__io_in_key_2_2),
    .io_in_key_2_3(xor__io_in_key_2_3),
    .io_in_key_3_0(xor__io_in_key_3_0),
    .io_in_key_3_1(xor__io_in_key_3_1),
    .io_in_key_3_2(xor__io_in_key_3_2),
    .io_in_key_3_3(xor__io_in_key_3_3)
  );
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 174:19]
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_XOR invxor ( // @[AES_PipelinedElasticBuffer.scala 184:22]
    .io_out_state_0_0(invxor_io_out_state_0_0),
    .io_out_state_0_1(invxor_io_out_state_0_1),
    .io_out_state_0_2(invxor_io_out_state_0_2),
    .io_out_state_0_3(invxor_io_out_state_0_3),
    .io_out_state_1_0(invxor_io_out_state_1_0),
    .io_out_state_1_1(invxor_io_out_state_1_1),
    .io_out_state_1_2(invxor_io_out_state_1_2),
    .io_out_state_1_3(invxor_io_out_state_1_3),
    .io_out_state_2_0(invxor_io_out_state_2_0),
    .io_out_state_2_1(invxor_io_out_state_2_1),
    .io_out_state_2_2(invxor_io_out_state_2_2),
    .io_out_state_2_3(invxor_io_out_state_2_3),
    .io_out_state_3_0(invxor_io_out_state_3_0),
    .io_out_state_3_1(invxor_io_out_state_3_1),
    .io_out_state_3_2(invxor_io_out_state_3_2),
    .io_out_state_3_3(invxor_io_out_state_3_3),
    .io_in_state_0_0(invxor_io_in_state_0_0),
    .io_in_state_0_1(invxor_io_in_state_0_1),
    .io_in_state_0_2(invxor_io_in_state_0_2),
    .io_in_state_0_3(invxor_io_in_state_0_3),
    .io_in_state_1_0(invxor_io_in_state_1_0),
    .io_in_state_1_1(invxor_io_in_state_1_1),
    .io_in_state_1_2(invxor_io_in_state_1_2),
    .io_in_state_1_3(invxor_io_in_state_1_3),
    .io_in_state_2_0(invxor_io_in_state_2_0),
    .io_in_state_2_1(invxor_io_in_state_2_1),
    .io_in_state_2_2(invxor_io_in_state_2_2),
    .io_in_state_2_3(invxor_io_in_state_2_3),
    .io_in_state_3_0(invxor_io_in_state_3_0),
    .io_in_state_3_1(invxor_io_in_state_3_1),
    .io_in_state_3_2(invxor_io_in_state_3_2),
    .io_in_state_3_3(invxor_io_in_state_3_3),
    .io_in_key_0_0(invxor_io_in_key_0_0),
    .io_in_key_0_1(invxor_io_in_key_0_1),
    .io_in_key_0_2(invxor_io_in_key_0_2),
    .io_in_key_0_3(invxor_io_in_key_0_3),
    .io_in_key_1_0(invxor_io_in_key_1_0),
    .io_in_key_1_1(invxor_io_in_key_1_1),
    .io_in_key_1_2(invxor_io_in_key_1_2),
    .io_in_key_1_3(invxor_io_in_key_1_3),
    .io_in_key_2_0(invxor_io_in_key_2_0),
    .io_in_key_2_1(invxor_io_in_key_2_1),
    .io_in_key_2_2(invxor_io_in_key_2_2),
    .io_in_key_2_3(invxor_io_in_key_2_3),
    .io_in_key_3_0(invxor_io_in_key_3_0),
    .io_in_key_3_1(invxor_io_in_key_3_1),
    .io_in_key_3_2(invxor_io_in_key_3_2),
    .io_in_key_3_3(invxor_io_in_key_3_3)
  );
  AES_InvMixColumns invmix ( // @[AES_PipelinedElasticBuffer.scala 189:22]
    .io_out_state_0_0(invmix_io_out_state_0_0),
    .io_out_state_0_1(invmix_io_out_state_0_1),
    .io_out_state_0_2(invmix_io_out_state_0_2),
    .io_out_state_0_3(invmix_io_out_state_0_3),
    .io_out_state_1_0(invmix_io_out_state_1_0),
    .io_out_state_1_1(invmix_io_out_state_1_1),
    .io_out_state_1_2(invmix_io_out_state_1_2),
    .io_out_state_1_3(invmix_io_out_state_1_3),
    .io_out_state_2_0(invmix_io_out_state_2_0),
    .io_out_state_2_1(invmix_io_out_state_2_1),
    .io_out_state_2_2(invmix_io_out_state_2_2),
    .io_out_state_2_3(invmix_io_out_state_2_3),
    .io_out_state_3_0(invmix_io_out_state_3_0),
    .io_out_state_3_1(invmix_io_out_state_3_1),
    .io_out_state_3_2(invmix_io_out_state_3_2),
    .io_out_state_3_3(invmix_io_out_state_3_3),
    .io_in_state_0_0(invmix_io_in_state_0_0),
    .io_in_state_0_1(invmix_io_in_state_0_1),
    .io_in_state_0_2(invmix_io_in_state_0_2),
    .io_in_state_0_3(invmix_io_in_state_0_3),
    .io_in_state_1_0(invmix_io_in_state_1_0),
    .io_in_state_1_1(invmix_io_in_state_1_1),
    .io_in_state_1_2(invmix_io_in_state_1_2),
    .io_in_state_1_3(invmix_io_in_state_1_3),
    .io_in_state_2_0(invmix_io_in_state_2_0),
    .io_in_state_2_1(invmix_io_in_state_2_1),
    .io_in_state_2_2(invmix_io_in_state_2_2),
    .io_in_state_2_3(invmix_io_in_state_2_3),
    .io_in_state_3_0(invmix_io_in_state_3_0),
    .io_in_state_3_1(invmix_io_in_state_3_1),
    .io_in_state_3_2(invmix_io_in_state_3_2),
    .io_in_state_3_3(invmix_io_in_state_3_3)
  );
  AES_InvShiftRows invshift ( // @[AES_PipelinedElasticBuffer.scala 192:24]
    .io_out_state_0_0(invshift_io_out_state_0_0),
    .io_out_state_0_1(invshift_io_out_state_0_1),
    .io_out_state_0_2(invshift_io_out_state_0_2),
    .io_out_state_0_3(invshift_io_out_state_0_3),
    .io_out_state_1_0(invshift_io_out_state_1_0),
    .io_out_state_1_1(invshift_io_out_state_1_1),
    .io_out_state_1_2(invshift_io_out_state_1_2),
    .io_out_state_1_3(invshift_io_out_state_1_3),
    .io_out_state_2_0(invshift_io_out_state_2_0),
    .io_out_state_2_1(invshift_io_out_state_2_1),
    .io_out_state_2_2(invshift_io_out_state_2_2),
    .io_out_state_2_3(invshift_io_out_state_2_3),
    .io_out_state_3_0(invshift_io_out_state_3_0),
    .io_out_state_3_1(invshift_io_out_state_3_1),
    .io_out_state_3_2(invshift_io_out_state_3_2),
    .io_out_state_3_3(invshift_io_out_state_3_3),
    .io_in_state_0_0(invshift_io_in_state_0_0),
    .io_in_state_0_1(invshift_io_in_state_0_1),
    .io_in_state_0_2(invshift_io_in_state_0_2),
    .io_in_state_0_3(invshift_io_in_state_0_3),
    .io_in_state_1_0(invshift_io_in_state_1_0),
    .io_in_state_1_1(invshift_io_in_state_1_1),
    .io_in_state_1_2(invshift_io_in_state_1_2),
    .io_in_state_1_3(invshift_io_in_state_1_3),
    .io_in_state_2_0(invshift_io_in_state_2_0),
    .io_in_state_2_1(invshift_io_in_state_2_1),
    .io_in_state_2_2(invshift_io_in_state_2_2),
    .io_in_state_2_3(invshift_io_in_state_2_3),
    .io_in_state_3_0(invshift_io_in_state_3_0),
    .io_in_state_3_1(invshift_io_in_state_3_1),
    .io_in_state_3_2(invshift_io_in_state_3_2),
    .io_in_state_3_3(invshift_io_in_state_3_3)
  );
  AES_InvSubBytes invsub ( // @[AES_PipelinedElasticBuffer.scala 199:22]
    .io_out_state_0_0(invsub_io_out_state_0_0),
    .io_out_state_0_1(invsub_io_out_state_0_1),
    .io_out_state_0_2(invsub_io_out_state_0_2),
    .io_out_state_0_3(invsub_io_out_state_0_3),
    .io_out_state_1_0(invsub_io_out_state_1_0),
    .io_out_state_1_1(invsub_io_out_state_1_1),
    .io_out_state_1_2(invsub_io_out_state_1_2),
    .io_out_state_1_3(invsub_io_out_state_1_3),
    .io_out_state_2_0(invsub_io_out_state_2_0),
    .io_out_state_2_1(invsub_io_out_state_2_1),
    .io_out_state_2_2(invsub_io_out_state_2_2),
    .io_out_state_2_3(invsub_io_out_state_2_3),
    .io_out_state_3_0(invsub_io_out_state_3_0),
    .io_out_state_3_1(invsub_io_out_state_3_1),
    .io_out_state_3_2(invsub_io_out_state_3_2),
    .io_out_state_3_3(invsub_io_out_state_3_3),
    .io_in_state_0_0(invsub_io_in_state_0_0),
    .io_in_state_0_1(invsub_io_in_state_0_1),
    .io_in_state_0_2(invsub_io_in_state_0_2),
    .io_in_state_0_3(invsub_io_in_state_0_3),
    .io_in_state_1_0(invsub_io_in_state_1_0),
    .io_in_state_1_1(invsub_io_in_state_1_1),
    .io_in_state_1_2(invsub_io_in_state_1_2),
    .io_in_state_1_3(invsub_io_in_state_1_3),
    .io_in_state_2_0(invsub_io_in_state_2_0),
    .io_in_state_2_1(invsub_io_in_state_2_1),
    .io_in_state_2_2(invsub_io_in_state_2_2),
    .io_in_state_2_3(invsub_io_in_state_2_3),
    .io_in_state_3_0(invsub_io_in_state_3_0),
    .io_in_state_3_1(invsub_io_in_state_3_1),
    .io_in_state_3_2(invsub_io_in_state_3_2),
    .io_in_state_3_3(invsub_io_in_state_3_3)
  );
  AES_GetNewKey_5 key ( // @[AES_PipelinedElasticBuffer.scala 202:19]
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  AES_InvGetNewKey_5 invkey ( // @[AES_PipelinedElasticBuffer.scala 206:22]
    .io_out_key_0_0(invkey_io_out_key_0_0),
    .io_out_key_0_1(invkey_io_out_key_0_1),
    .io_out_key_0_2(invkey_io_out_key_0_2),
    .io_out_key_0_3(invkey_io_out_key_0_3),
    .io_out_key_1_0(invkey_io_out_key_1_0),
    .io_out_key_1_1(invkey_io_out_key_1_1),
    .io_out_key_1_2(invkey_io_out_key_1_2),
    .io_out_key_1_3(invkey_io_out_key_1_3),
    .io_out_key_2_0(invkey_io_out_key_2_0),
    .io_out_key_2_1(invkey_io_out_key_2_1),
    .io_out_key_2_2(invkey_io_out_key_2_2),
    .io_out_key_2_3(invkey_io_out_key_2_3),
    .io_out_key_3_0(invkey_io_out_key_3_0),
    .io_out_key_3_1(invkey_io_out_key_3_1),
    .io_out_key_3_2(invkey_io_out_key_3_2),
    .io_out_key_3_3(invkey_io_out_key_3_3),
    .io_in_key_0_0(invkey_io_in_key_0_0),
    .io_in_key_0_1(invkey_io_in_key_0_1),
    .io_in_key_0_2(invkey_io_in_key_0_2),
    .io_in_key_0_3(invkey_io_in_key_0_3),
    .io_in_key_1_0(invkey_io_in_key_1_0),
    .io_in_key_1_1(invkey_io_in_key_1_1),
    .io_in_key_1_2(invkey_io_in_key_1_2),
    .io_in_key_1_3(invkey_io_in_key_1_3),
    .io_in_key_2_0(invkey_io_in_key_2_0),
    .io_in_key_2_1(invkey_io_in_key_2_1),
    .io_in_key_2_2(invkey_io_in_key_2_2),
    .io_in_key_2_3(invkey_io_in_key_2_3),
    .io_in_key_3_0(invkey_io_in_key_3_0),
    .io_in_key_3_1(invkey_io_in_key_3_1),
    .io_in_key_3_2(invkey_io_in_key_3_2),
    .io_in_key_3_3(invkey_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 151:27]
  assign io_out_bits_state_0_0 = invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_1 = invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_2 = invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_3 = invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_0 = invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_1 = invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_2 = invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_3 = invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_0 = invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_1 = invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_2 = invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_3 = invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_0 = invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_1 = invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_2 = invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_3 = invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_0 = invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_1 = invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_2 = invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_3 = invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_0 = invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_1 = invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_2 = invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_3 = invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_0 = invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_1 = invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_2 = invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_3 = invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_0 = invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_1 = invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_2 = invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_3 = invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 150:18]
  assign xor__io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign sub_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign invxor_io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invmix_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invshift_io_in_state_0_0 = invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_1 = invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_2 = invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_3 = invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_0 = invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_1 = invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_2 = invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_3 = invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_0 = invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_1 = invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_2 = invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_3 = invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_0 = invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_1 = invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_2 = invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_3 = invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invsub_io_in_state_0_0 = invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_1 = invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_2 = invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_3 = invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_0 = invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_1 = invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_2 = invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_3 = invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_0 = invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_1 = invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_2 = invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_3 = invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_0 = invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_1 = invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_2 = invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_3 = invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 146:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 146:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 165:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 159:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_6(
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 237:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 240:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 241:13]
endmodule
module AES_InvGetNewKey_6(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] w4 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w5 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w6 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [31:0] w7 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] w3 = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  wire [31:0] w2 = w6 ^ w5; // @[AES_PipelinedElasticBuffer.scala 301:12]
  wire [31:0] w1 = w5 ^ w4; // @[AES_PipelinedElasticBuffer.scala 302:12]
  wire [31:0] temp = 32'h8000000 ^ sub_io_out; // @[AES_PipelinedElasticBuffer.scala 310:16]
  wire [31:0] w0 = w4 ^ temp; // @[AES_PipelinedElasticBuffer.scala 303:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 305:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 308:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w0[31:24]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_1 = w0[23:16]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_2 = w0[15:8]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_3 = w0[7:0]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_1_0 = w1[31:24]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_1 = w1[23:16]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_2 = w1[15:8]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_3 = w1[7:0]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_2_0 = w2[31:24]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_1 = w2[23:16]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_2 = w2[15:8]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_3 = w2[7:0]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_3_0 = w3[31:24]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_1 = w3[23:16]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_2 = w3[15:8]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_3 = w3[7:0]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign rot_io_in = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 309:13]
endmodule
module AES_ProcessingElement_6(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 146:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:23 AES_PipelinedElasticBuffer.scala 156:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 163:21 AES_PipelinedElasticBuffer.scala 163:21]
  AES_XOR xor_ ( // @[AES_PipelinedElasticBuffer.scala 169:19]
    .io_out_state_0_0(xor__io_out_state_0_0),
    .io_out_state_0_1(xor__io_out_state_0_1),
    .io_out_state_0_2(xor__io_out_state_0_2),
    .io_out_state_0_3(xor__io_out_state_0_3),
    .io_out_state_1_0(xor__io_out_state_1_0),
    .io_out_state_1_1(xor__io_out_state_1_1),
    .io_out_state_1_2(xor__io_out_state_1_2),
    .io_out_state_1_3(xor__io_out_state_1_3),
    .io_out_state_2_0(xor__io_out_state_2_0),
    .io_out_state_2_1(xor__io_out_state_2_1),
    .io_out_state_2_2(xor__io_out_state_2_2),
    .io_out_state_2_3(xor__io_out_state_2_3),
    .io_out_state_3_0(xor__io_out_state_3_0),
    .io_out_state_3_1(xor__io_out_state_3_1),
    .io_out_state_3_2(xor__io_out_state_3_2),
    .io_out_state_3_3(xor__io_out_state_3_3),
    .io_in_state_0_0(xor__io_in_state_0_0),
    .io_in_state_0_1(xor__io_in_state_0_1),
    .io_in_state_0_2(xor__io_in_state_0_2),
    .io_in_state_0_3(xor__io_in_state_0_3),
    .io_in_state_1_0(xor__io_in_state_1_0),
    .io_in_state_1_1(xor__io_in_state_1_1),
    .io_in_state_1_2(xor__io_in_state_1_2),
    .io_in_state_1_3(xor__io_in_state_1_3),
    .io_in_state_2_0(xor__io_in_state_2_0),
    .io_in_state_2_1(xor__io_in_state_2_1),
    .io_in_state_2_2(xor__io_in_state_2_2),
    .io_in_state_2_3(xor__io_in_state_2_3),
    .io_in_state_3_0(xor__io_in_state_3_0),
    .io_in_state_3_1(xor__io_in_state_3_1),
    .io_in_state_3_2(xor__io_in_state_3_2),
    .io_in_state_3_3(xor__io_in_state_3_3),
    .io_in_key_0_0(xor__io_in_key_0_0),
    .io_in_key_0_1(xor__io_in_key_0_1),
    .io_in_key_0_2(xor__io_in_key_0_2),
    .io_in_key_0_3(xor__io_in_key_0_3),
    .io_in_key_1_0(xor__io_in_key_1_0),
    .io_in_key_1_1(xor__io_in_key_1_1),
    .io_in_key_1_2(xor__io_in_key_1_2),
    .io_in_key_1_3(xor__io_in_key_1_3),
    .io_in_key_2_0(xor__io_in_key_2_0),
    .io_in_key_2_1(xor__io_in_key_2_1),
    .io_in_key_2_2(xor__io_in_key_2_2),
    .io_in_key_2_3(xor__io_in_key_2_3),
    .io_in_key_3_0(xor__io_in_key_3_0),
    .io_in_key_3_1(xor__io_in_key_3_1),
    .io_in_key_3_2(xor__io_in_key_3_2),
    .io_in_key_3_3(xor__io_in_key_3_3)
  );
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 174:19]
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_XOR invxor ( // @[AES_PipelinedElasticBuffer.scala 184:22]
    .io_out_state_0_0(invxor_io_out_state_0_0),
    .io_out_state_0_1(invxor_io_out_state_0_1),
    .io_out_state_0_2(invxor_io_out_state_0_2),
    .io_out_state_0_3(invxor_io_out_state_0_3),
    .io_out_state_1_0(invxor_io_out_state_1_0),
    .io_out_state_1_1(invxor_io_out_state_1_1),
    .io_out_state_1_2(invxor_io_out_state_1_2),
    .io_out_state_1_3(invxor_io_out_state_1_3),
    .io_out_state_2_0(invxor_io_out_state_2_0),
    .io_out_state_2_1(invxor_io_out_state_2_1),
    .io_out_state_2_2(invxor_io_out_state_2_2),
    .io_out_state_2_3(invxor_io_out_state_2_3),
    .io_out_state_3_0(invxor_io_out_state_3_0),
    .io_out_state_3_1(invxor_io_out_state_3_1),
    .io_out_state_3_2(invxor_io_out_state_3_2),
    .io_out_state_3_3(invxor_io_out_state_3_3),
    .io_in_state_0_0(invxor_io_in_state_0_0),
    .io_in_state_0_1(invxor_io_in_state_0_1),
    .io_in_state_0_2(invxor_io_in_state_0_2),
    .io_in_state_0_3(invxor_io_in_state_0_3),
    .io_in_state_1_0(invxor_io_in_state_1_0),
    .io_in_state_1_1(invxor_io_in_state_1_1),
    .io_in_state_1_2(invxor_io_in_state_1_2),
    .io_in_state_1_3(invxor_io_in_state_1_3),
    .io_in_state_2_0(invxor_io_in_state_2_0),
    .io_in_state_2_1(invxor_io_in_state_2_1),
    .io_in_state_2_2(invxor_io_in_state_2_2),
    .io_in_state_2_3(invxor_io_in_state_2_3),
    .io_in_state_3_0(invxor_io_in_state_3_0),
    .io_in_state_3_1(invxor_io_in_state_3_1),
    .io_in_state_3_2(invxor_io_in_state_3_2),
    .io_in_state_3_3(invxor_io_in_state_3_3),
    .io_in_key_0_0(invxor_io_in_key_0_0),
    .io_in_key_0_1(invxor_io_in_key_0_1),
    .io_in_key_0_2(invxor_io_in_key_0_2),
    .io_in_key_0_3(invxor_io_in_key_0_3),
    .io_in_key_1_0(invxor_io_in_key_1_0),
    .io_in_key_1_1(invxor_io_in_key_1_1),
    .io_in_key_1_2(invxor_io_in_key_1_2),
    .io_in_key_1_3(invxor_io_in_key_1_3),
    .io_in_key_2_0(invxor_io_in_key_2_0),
    .io_in_key_2_1(invxor_io_in_key_2_1),
    .io_in_key_2_2(invxor_io_in_key_2_2),
    .io_in_key_2_3(invxor_io_in_key_2_3),
    .io_in_key_3_0(invxor_io_in_key_3_0),
    .io_in_key_3_1(invxor_io_in_key_3_1),
    .io_in_key_3_2(invxor_io_in_key_3_2),
    .io_in_key_3_3(invxor_io_in_key_3_3)
  );
  AES_InvMixColumns invmix ( // @[AES_PipelinedElasticBuffer.scala 189:22]
    .io_out_state_0_0(invmix_io_out_state_0_0),
    .io_out_state_0_1(invmix_io_out_state_0_1),
    .io_out_state_0_2(invmix_io_out_state_0_2),
    .io_out_state_0_3(invmix_io_out_state_0_3),
    .io_out_state_1_0(invmix_io_out_state_1_0),
    .io_out_state_1_1(invmix_io_out_state_1_1),
    .io_out_state_1_2(invmix_io_out_state_1_2),
    .io_out_state_1_3(invmix_io_out_state_1_3),
    .io_out_state_2_0(invmix_io_out_state_2_0),
    .io_out_state_2_1(invmix_io_out_state_2_1),
    .io_out_state_2_2(invmix_io_out_state_2_2),
    .io_out_state_2_3(invmix_io_out_state_2_3),
    .io_out_state_3_0(invmix_io_out_state_3_0),
    .io_out_state_3_1(invmix_io_out_state_3_1),
    .io_out_state_3_2(invmix_io_out_state_3_2),
    .io_out_state_3_3(invmix_io_out_state_3_3),
    .io_in_state_0_0(invmix_io_in_state_0_0),
    .io_in_state_0_1(invmix_io_in_state_0_1),
    .io_in_state_0_2(invmix_io_in_state_0_2),
    .io_in_state_0_3(invmix_io_in_state_0_3),
    .io_in_state_1_0(invmix_io_in_state_1_0),
    .io_in_state_1_1(invmix_io_in_state_1_1),
    .io_in_state_1_2(invmix_io_in_state_1_2),
    .io_in_state_1_3(invmix_io_in_state_1_3),
    .io_in_state_2_0(invmix_io_in_state_2_0),
    .io_in_state_2_1(invmix_io_in_state_2_1),
    .io_in_state_2_2(invmix_io_in_state_2_2),
    .io_in_state_2_3(invmix_io_in_state_2_3),
    .io_in_state_3_0(invmix_io_in_state_3_0),
    .io_in_state_3_1(invmix_io_in_state_3_1),
    .io_in_state_3_2(invmix_io_in_state_3_2),
    .io_in_state_3_3(invmix_io_in_state_3_3)
  );
  AES_InvShiftRows invshift ( // @[AES_PipelinedElasticBuffer.scala 192:24]
    .io_out_state_0_0(invshift_io_out_state_0_0),
    .io_out_state_0_1(invshift_io_out_state_0_1),
    .io_out_state_0_2(invshift_io_out_state_0_2),
    .io_out_state_0_3(invshift_io_out_state_0_3),
    .io_out_state_1_0(invshift_io_out_state_1_0),
    .io_out_state_1_1(invshift_io_out_state_1_1),
    .io_out_state_1_2(invshift_io_out_state_1_2),
    .io_out_state_1_3(invshift_io_out_state_1_3),
    .io_out_state_2_0(invshift_io_out_state_2_0),
    .io_out_state_2_1(invshift_io_out_state_2_1),
    .io_out_state_2_2(invshift_io_out_state_2_2),
    .io_out_state_2_3(invshift_io_out_state_2_3),
    .io_out_state_3_0(invshift_io_out_state_3_0),
    .io_out_state_3_1(invshift_io_out_state_3_1),
    .io_out_state_3_2(invshift_io_out_state_3_2),
    .io_out_state_3_3(invshift_io_out_state_3_3),
    .io_in_state_0_0(invshift_io_in_state_0_0),
    .io_in_state_0_1(invshift_io_in_state_0_1),
    .io_in_state_0_2(invshift_io_in_state_0_2),
    .io_in_state_0_3(invshift_io_in_state_0_3),
    .io_in_state_1_0(invshift_io_in_state_1_0),
    .io_in_state_1_1(invshift_io_in_state_1_1),
    .io_in_state_1_2(invshift_io_in_state_1_2),
    .io_in_state_1_3(invshift_io_in_state_1_3),
    .io_in_state_2_0(invshift_io_in_state_2_0),
    .io_in_state_2_1(invshift_io_in_state_2_1),
    .io_in_state_2_2(invshift_io_in_state_2_2),
    .io_in_state_2_3(invshift_io_in_state_2_3),
    .io_in_state_3_0(invshift_io_in_state_3_0),
    .io_in_state_3_1(invshift_io_in_state_3_1),
    .io_in_state_3_2(invshift_io_in_state_3_2),
    .io_in_state_3_3(invshift_io_in_state_3_3)
  );
  AES_InvSubBytes invsub ( // @[AES_PipelinedElasticBuffer.scala 199:22]
    .io_out_state_0_0(invsub_io_out_state_0_0),
    .io_out_state_0_1(invsub_io_out_state_0_1),
    .io_out_state_0_2(invsub_io_out_state_0_2),
    .io_out_state_0_3(invsub_io_out_state_0_3),
    .io_out_state_1_0(invsub_io_out_state_1_0),
    .io_out_state_1_1(invsub_io_out_state_1_1),
    .io_out_state_1_2(invsub_io_out_state_1_2),
    .io_out_state_1_3(invsub_io_out_state_1_3),
    .io_out_state_2_0(invsub_io_out_state_2_0),
    .io_out_state_2_1(invsub_io_out_state_2_1),
    .io_out_state_2_2(invsub_io_out_state_2_2),
    .io_out_state_2_3(invsub_io_out_state_2_3),
    .io_out_state_3_0(invsub_io_out_state_3_0),
    .io_out_state_3_1(invsub_io_out_state_3_1),
    .io_out_state_3_2(invsub_io_out_state_3_2),
    .io_out_state_3_3(invsub_io_out_state_3_3),
    .io_in_state_0_0(invsub_io_in_state_0_0),
    .io_in_state_0_1(invsub_io_in_state_0_1),
    .io_in_state_0_2(invsub_io_in_state_0_2),
    .io_in_state_0_3(invsub_io_in_state_0_3),
    .io_in_state_1_0(invsub_io_in_state_1_0),
    .io_in_state_1_1(invsub_io_in_state_1_1),
    .io_in_state_1_2(invsub_io_in_state_1_2),
    .io_in_state_1_3(invsub_io_in_state_1_3),
    .io_in_state_2_0(invsub_io_in_state_2_0),
    .io_in_state_2_1(invsub_io_in_state_2_1),
    .io_in_state_2_2(invsub_io_in_state_2_2),
    .io_in_state_2_3(invsub_io_in_state_2_3),
    .io_in_state_3_0(invsub_io_in_state_3_0),
    .io_in_state_3_1(invsub_io_in_state_3_1),
    .io_in_state_3_2(invsub_io_in_state_3_2),
    .io_in_state_3_3(invsub_io_in_state_3_3)
  );
  AES_GetNewKey_6 key ( // @[AES_PipelinedElasticBuffer.scala 202:19]
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  AES_InvGetNewKey_6 invkey ( // @[AES_PipelinedElasticBuffer.scala 206:22]
    .io_out_key_0_0(invkey_io_out_key_0_0),
    .io_out_key_0_1(invkey_io_out_key_0_1),
    .io_out_key_0_2(invkey_io_out_key_0_2),
    .io_out_key_0_3(invkey_io_out_key_0_3),
    .io_out_key_1_0(invkey_io_out_key_1_0),
    .io_out_key_1_1(invkey_io_out_key_1_1),
    .io_out_key_1_2(invkey_io_out_key_1_2),
    .io_out_key_1_3(invkey_io_out_key_1_3),
    .io_out_key_2_0(invkey_io_out_key_2_0),
    .io_out_key_2_1(invkey_io_out_key_2_1),
    .io_out_key_2_2(invkey_io_out_key_2_2),
    .io_out_key_2_3(invkey_io_out_key_2_3),
    .io_out_key_3_0(invkey_io_out_key_3_0),
    .io_out_key_3_1(invkey_io_out_key_3_1),
    .io_out_key_3_2(invkey_io_out_key_3_2),
    .io_out_key_3_3(invkey_io_out_key_3_3),
    .io_in_key_0_0(invkey_io_in_key_0_0),
    .io_in_key_0_1(invkey_io_in_key_0_1),
    .io_in_key_0_2(invkey_io_in_key_0_2),
    .io_in_key_0_3(invkey_io_in_key_0_3),
    .io_in_key_1_0(invkey_io_in_key_1_0),
    .io_in_key_1_1(invkey_io_in_key_1_1),
    .io_in_key_1_2(invkey_io_in_key_1_2),
    .io_in_key_1_3(invkey_io_in_key_1_3),
    .io_in_key_2_0(invkey_io_in_key_2_0),
    .io_in_key_2_1(invkey_io_in_key_2_1),
    .io_in_key_2_2(invkey_io_in_key_2_2),
    .io_in_key_2_3(invkey_io_in_key_2_3),
    .io_in_key_3_0(invkey_io_in_key_3_0),
    .io_in_key_3_1(invkey_io_in_key_3_1),
    .io_in_key_3_2(invkey_io_in_key_3_2),
    .io_in_key_3_3(invkey_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 151:27]
  assign io_out_bits_state_0_0 = invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_1 = invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_2 = invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_3 = invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_0 = invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_1 = invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_2 = invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_3 = invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_0 = invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_1 = invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_2 = invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_3 = invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_0 = invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_1 = invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_2 = invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_3 = invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_0 = invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_1 = invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_2 = invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_3 = invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_0 = invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_1 = invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_2 = invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_3 = invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_0 = invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_1 = invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_2 = invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_3 = invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_0 = invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_1 = invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_2 = invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_3 = invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 150:18]
  assign xor__io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign sub_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign invxor_io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invmix_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invshift_io_in_state_0_0 = invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_1 = invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_2 = invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_3 = invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_0 = invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_1 = invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_2 = invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_3 = invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_0 = invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_1 = invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_2 = invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_3 = invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_0 = invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_1 = invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_2 = invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_3 = invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invsub_io_in_state_0_0 = invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_1 = invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_2 = invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_3 = invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_0 = invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_1 = invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_2 = invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_3 = invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_0 = invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_1 = invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_2 = invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_3 = invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_0 = invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_1 = invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_2 = invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_3 = invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 146:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 146:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 165:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 159:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_7(
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 237:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 240:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 241:13]
endmodule
module AES_InvGetNewKey_7(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] w4 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w5 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w6 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [31:0] w7 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] w3 = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  wire [31:0] w2 = w6 ^ w5; // @[AES_PipelinedElasticBuffer.scala 301:12]
  wire [31:0] w1 = w5 ^ w4; // @[AES_PipelinedElasticBuffer.scala 302:12]
  wire [31:0] temp = 32'h4000000 ^ sub_io_out; // @[AES_PipelinedElasticBuffer.scala 310:16]
  wire [31:0] w0 = w4 ^ temp; // @[AES_PipelinedElasticBuffer.scala 303:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 305:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 308:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w0[31:24]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_1 = w0[23:16]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_2 = w0[15:8]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_3 = w0[7:0]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_1_0 = w1[31:24]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_1 = w1[23:16]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_2 = w1[15:8]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_3 = w1[7:0]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_2_0 = w2[31:24]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_1 = w2[23:16]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_2 = w2[15:8]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_3 = w2[7:0]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_3_0 = w3[31:24]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_1 = w3[23:16]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_2 = w3[15:8]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_3 = w3[7:0]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign rot_io_in = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 309:13]
endmodule
module AES_ProcessingElement_7(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 146:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:23 AES_PipelinedElasticBuffer.scala 156:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 163:21 AES_PipelinedElasticBuffer.scala 163:21]
  AES_XOR xor_ ( // @[AES_PipelinedElasticBuffer.scala 169:19]
    .io_out_state_0_0(xor__io_out_state_0_0),
    .io_out_state_0_1(xor__io_out_state_0_1),
    .io_out_state_0_2(xor__io_out_state_0_2),
    .io_out_state_0_3(xor__io_out_state_0_3),
    .io_out_state_1_0(xor__io_out_state_1_0),
    .io_out_state_1_1(xor__io_out_state_1_1),
    .io_out_state_1_2(xor__io_out_state_1_2),
    .io_out_state_1_3(xor__io_out_state_1_3),
    .io_out_state_2_0(xor__io_out_state_2_0),
    .io_out_state_2_1(xor__io_out_state_2_1),
    .io_out_state_2_2(xor__io_out_state_2_2),
    .io_out_state_2_3(xor__io_out_state_2_3),
    .io_out_state_3_0(xor__io_out_state_3_0),
    .io_out_state_3_1(xor__io_out_state_3_1),
    .io_out_state_3_2(xor__io_out_state_3_2),
    .io_out_state_3_3(xor__io_out_state_3_3),
    .io_in_state_0_0(xor__io_in_state_0_0),
    .io_in_state_0_1(xor__io_in_state_0_1),
    .io_in_state_0_2(xor__io_in_state_0_2),
    .io_in_state_0_3(xor__io_in_state_0_3),
    .io_in_state_1_0(xor__io_in_state_1_0),
    .io_in_state_1_1(xor__io_in_state_1_1),
    .io_in_state_1_2(xor__io_in_state_1_2),
    .io_in_state_1_3(xor__io_in_state_1_3),
    .io_in_state_2_0(xor__io_in_state_2_0),
    .io_in_state_2_1(xor__io_in_state_2_1),
    .io_in_state_2_2(xor__io_in_state_2_2),
    .io_in_state_2_3(xor__io_in_state_2_3),
    .io_in_state_3_0(xor__io_in_state_3_0),
    .io_in_state_3_1(xor__io_in_state_3_1),
    .io_in_state_3_2(xor__io_in_state_3_2),
    .io_in_state_3_3(xor__io_in_state_3_3),
    .io_in_key_0_0(xor__io_in_key_0_0),
    .io_in_key_0_1(xor__io_in_key_0_1),
    .io_in_key_0_2(xor__io_in_key_0_2),
    .io_in_key_0_3(xor__io_in_key_0_3),
    .io_in_key_1_0(xor__io_in_key_1_0),
    .io_in_key_1_1(xor__io_in_key_1_1),
    .io_in_key_1_2(xor__io_in_key_1_2),
    .io_in_key_1_3(xor__io_in_key_1_3),
    .io_in_key_2_0(xor__io_in_key_2_0),
    .io_in_key_2_1(xor__io_in_key_2_1),
    .io_in_key_2_2(xor__io_in_key_2_2),
    .io_in_key_2_3(xor__io_in_key_2_3),
    .io_in_key_3_0(xor__io_in_key_3_0),
    .io_in_key_3_1(xor__io_in_key_3_1),
    .io_in_key_3_2(xor__io_in_key_3_2),
    .io_in_key_3_3(xor__io_in_key_3_3)
  );
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 174:19]
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_XOR invxor ( // @[AES_PipelinedElasticBuffer.scala 184:22]
    .io_out_state_0_0(invxor_io_out_state_0_0),
    .io_out_state_0_1(invxor_io_out_state_0_1),
    .io_out_state_0_2(invxor_io_out_state_0_2),
    .io_out_state_0_3(invxor_io_out_state_0_3),
    .io_out_state_1_0(invxor_io_out_state_1_0),
    .io_out_state_1_1(invxor_io_out_state_1_1),
    .io_out_state_1_2(invxor_io_out_state_1_2),
    .io_out_state_1_3(invxor_io_out_state_1_3),
    .io_out_state_2_0(invxor_io_out_state_2_0),
    .io_out_state_2_1(invxor_io_out_state_2_1),
    .io_out_state_2_2(invxor_io_out_state_2_2),
    .io_out_state_2_3(invxor_io_out_state_2_3),
    .io_out_state_3_0(invxor_io_out_state_3_0),
    .io_out_state_3_1(invxor_io_out_state_3_1),
    .io_out_state_3_2(invxor_io_out_state_3_2),
    .io_out_state_3_3(invxor_io_out_state_3_3),
    .io_in_state_0_0(invxor_io_in_state_0_0),
    .io_in_state_0_1(invxor_io_in_state_0_1),
    .io_in_state_0_2(invxor_io_in_state_0_2),
    .io_in_state_0_3(invxor_io_in_state_0_3),
    .io_in_state_1_0(invxor_io_in_state_1_0),
    .io_in_state_1_1(invxor_io_in_state_1_1),
    .io_in_state_1_2(invxor_io_in_state_1_2),
    .io_in_state_1_3(invxor_io_in_state_1_3),
    .io_in_state_2_0(invxor_io_in_state_2_0),
    .io_in_state_2_1(invxor_io_in_state_2_1),
    .io_in_state_2_2(invxor_io_in_state_2_2),
    .io_in_state_2_3(invxor_io_in_state_2_3),
    .io_in_state_3_0(invxor_io_in_state_3_0),
    .io_in_state_3_1(invxor_io_in_state_3_1),
    .io_in_state_3_2(invxor_io_in_state_3_2),
    .io_in_state_3_3(invxor_io_in_state_3_3),
    .io_in_key_0_0(invxor_io_in_key_0_0),
    .io_in_key_0_1(invxor_io_in_key_0_1),
    .io_in_key_0_2(invxor_io_in_key_0_2),
    .io_in_key_0_3(invxor_io_in_key_0_3),
    .io_in_key_1_0(invxor_io_in_key_1_0),
    .io_in_key_1_1(invxor_io_in_key_1_1),
    .io_in_key_1_2(invxor_io_in_key_1_2),
    .io_in_key_1_3(invxor_io_in_key_1_3),
    .io_in_key_2_0(invxor_io_in_key_2_0),
    .io_in_key_2_1(invxor_io_in_key_2_1),
    .io_in_key_2_2(invxor_io_in_key_2_2),
    .io_in_key_2_3(invxor_io_in_key_2_3),
    .io_in_key_3_0(invxor_io_in_key_3_0),
    .io_in_key_3_1(invxor_io_in_key_3_1),
    .io_in_key_3_2(invxor_io_in_key_3_2),
    .io_in_key_3_3(invxor_io_in_key_3_3)
  );
  AES_InvMixColumns invmix ( // @[AES_PipelinedElasticBuffer.scala 189:22]
    .io_out_state_0_0(invmix_io_out_state_0_0),
    .io_out_state_0_1(invmix_io_out_state_0_1),
    .io_out_state_0_2(invmix_io_out_state_0_2),
    .io_out_state_0_3(invmix_io_out_state_0_3),
    .io_out_state_1_0(invmix_io_out_state_1_0),
    .io_out_state_1_1(invmix_io_out_state_1_1),
    .io_out_state_1_2(invmix_io_out_state_1_2),
    .io_out_state_1_3(invmix_io_out_state_1_3),
    .io_out_state_2_0(invmix_io_out_state_2_0),
    .io_out_state_2_1(invmix_io_out_state_2_1),
    .io_out_state_2_2(invmix_io_out_state_2_2),
    .io_out_state_2_3(invmix_io_out_state_2_3),
    .io_out_state_3_0(invmix_io_out_state_3_0),
    .io_out_state_3_1(invmix_io_out_state_3_1),
    .io_out_state_3_2(invmix_io_out_state_3_2),
    .io_out_state_3_3(invmix_io_out_state_3_3),
    .io_in_state_0_0(invmix_io_in_state_0_0),
    .io_in_state_0_1(invmix_io_in_state_0_1),
    .io_in_state_0_2(invmix_io_in_state_0_2),
    .io_in_state_0_3(invmix_io_in_state_0_3),
    .io_in_state_1_0(invmix_io_in_state_1_0),
    .io_in_state_1_1(invmix_io_in_state_1_1),
    .io_in_state_1_2(invmix_io_in_state_1_2),
    .io_in_state_1_3(invmix_io_in_state_1_3),
    .io_in_state_2_0(invmix_io_in_state_2_0),
    .io_in_state_2_1(invmix_io_in_state_2_1),
    .io_in_state_2_2(invmix_io_in_state_2_2),
    .io_in_state_2_3(invmix_io_in_state_2_3),
    .io_in_state_3_0(invmix_io_in_state_3_0),
    .io_in_state_3_1(invmix_io_in_state_3_1),
    .io_in_state_3_2(invmix_io_in_state_3_2),
    .io_in_state_3_3(invmix_io_in_state_3_3)
  );
  AES_InvShiftRows invshift ( // @[AES_PipelinedElasticBuffer.scala 192:24]
    .io_out_state_0_0(invshift_io_out_state_0_0),
    .io_out_state_0_1(invshift_io_out_state_0_1),
    .io_out_state_0_2(invshift_io_out_state_0_2),
    .io_out_state_0_3(invshift_io_out_state_0_3),
    .io_out_state_1_0(invshift_io_out_state_1_0),
    .io_out_state_1_1(invshift_io_out_state_1_1),
    .io_out_state_1_2(invshift_io_out_state_1_2),
    .io_out_state_1_3(invshift_io_out_state_1_3),
    .io_out_state_2_0(invshift_io_out_state_2_0),
    .io_out_state_2_1(invshift_io_out_state_2_1),
    .io_out_state_2_2(invshift_io_out_state_2_2),
    .io_out_state_2_3(invshift_io_out_state_2_3),
    .io_out_state_3_0(invshift_io_out_state_3_0),
    .io_out_state_3_1(invshift_io_out_state_3_1),
    .io_out_state_3_2(invshift_io_out_state_3_2),
    .io_out_state_3_3(invshift_io_out_state_3_3),
    .io_in_state_0_0(invshift_io_in_state_0_0),
    .io_in_state_0_1(invshift_io_in_state_0_1),
    .io_in_state_0_2(invshift_io_in_state_0_2),
    .io_in_state_0_3(invshift_io_in_state_0_3),
    .io_in_state_1_0(invshift_io_in_state_1_0),
    .io_in_state_1_1(invshift_io_in_state_1_1),
    .io_in_state_1_2(invshift_io_in_state_1_2),
    .io_in_state_1_3(invshift_io_in_state_1_3),
    .io_in_state_2_0(invshift_io_in_state_2_0),
    .io_in_state_2_1(invshift_io_in_state_2_1),
    .io_in_state_2_2(invshift_io_in_state_2_2),
    .io_in_state_2_3(invshift_io_in_state_2_3),
    .io_in_state_3_0(invshift_io_in_state_3_0),
    .io_in_state_3_1(invshift_io_in_state_3_1),
    .io_in_state_3_2(invshift_io_in_state_3_2),
    .io_in_state_3_3(invshift_io_in_state_3_3)
  );
  AES_InvSubBytes invsub ( // @[AES_PipelinedElasticBuffer.scala 199:22]
    .io_out_state_0_0(invsub_io_out_state_0_0),
    .io_out_state_0_1(invsub_io_out_state_0_1),
    .io_out_state_0_2(invsub_io_out_state_0_2),
    .io_out_state_0_3(invsub_io_out_state_0_3),
    .io_out_state_1_0(invsub_io_out_state_1_0),
    .io_out_state_1_1(invsub_io_out_state_1_1),
    .io_out_state_1_2(invsub_io_out_state_1_2),
    .io_out_state_1_3(invsub_io_out_state_1_3),
    .io_out_state_2_0(invsub_io_out_state_2_0),
    .io_out_state_2_1(invsub_io_out_state_2_1),
    .io_out_state_2_2(invsub_io_out_state_2_2),
    .io_out_state_2_3(invsub_io_out_state_2_3),
    .io_out_state_3_0(invsub_io_out_state_3_0),
    .io_out_state_3_1(invsub_io_out_state_3_1),
    .io_out_state_3_2(invsub_io_out_state_3_2),
    .io_out_state_3_3(invsub_io_out_state_3_3),
    .io_in_state_0_0(invsub_io_in_state_0_0),
    .io_in_state_0_1(invsub_io_in_state_0_1),
    .io_in_state_0_2(invsub_io_in_state_0_2),
    .io_in_state_0_3(invsub_io_in_state_0_3),
    .io_in_state_1_0(invsub_io_in_state_1_0),
    .io_in_state_1_1(invsub_io_in_state_1_1),
    .io_in_state_1_2(invsub_io_in_state_1_2),
    .io_in_state_1_3(invsub_io_in_state_1_3),
    .io_in_state_2_0(invsub_io_in_state_2_0),
    .io_in_state_2_1(invsub_io_in_state_2_1),
    .io_in_state_2_2(invsub_io_in_state_2_2),
    .io_in_state_2_3(invsub_io_in_state_2_3),
    .io_in_state_3_0(invsub_io_in_state_3_0),
    .io_in_state_3_1(invsub_io_in_state_3_1),
    .io_in_state_3_2(invsub_io_in_state_3_2),
    .io_in_state_3_3(invsub_io_in_state_3_3)
  );
  AES_GetNewKey_7 key ( // @[AES_PipelinedElasticBuffer.scala 202:19]
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  AES_InvGetNewKey_7 invkey ( // @[AES_PipelinedElasticBuffer.scala 206:22]
    .io_out_key_0_0(invkey_io_out_key_0_0),
    .io_out_key_0_1(invkey_io_out_key_0_1),
    .io_out_key_0_2(invkey_io_out_key_0_2),
    .io_out_key_0_3(invkey_io_out_key_0_3),
    .io_out_key_1_0(invkey_io_out_key_1_0),
    .io_out_key_1_1(invkey_io_out_key_1_1),
    .io_out_key_1_2(invkey_io_out_key_1_2),
    .io_out_key_1_3(invkey_io_out_key_1_3),
    .io_out_key_2_0(invkey_io_out_key_2_0),
    .io_out_key_2_1(invkey_io_out_key_2_1),
    .io_out_key_2_2(invkey_io_out_key_2_2),
    .io_out_key_2_3(invkey_io_out_key_2_3),
    .io_out_key_3_0(invkey_io_out_key_3_0),
    .io_out_key_3_1(invkey_io_out_key_3_1),
    .io_out_key_3_2(invkey_io_out_key_3_2),
    .io_out_key_3_3(invkey_io_out_key_3_3),
    .io_in_key_0_0(invkey_io_in_key_0_0),
    .io_in_key_0_1(invkey_io_in_key_0_1),
    .io_in_key_0_2(invkey_io_in_key_0_2),
    .io_in_key_0_3(invkey_io_in_key_0_3),
    .io_in_key_1_0(invkey_io_in_key_1_0),
    .io_in_key_1_1(invkey_io_in_key_1_1),
    .io_in_key_1_2(invkey_io_in_key_1_2),
    .io_in_key_1_3(invkey_io_in_key_1_3),
    .io_in_key_2_0(invkey_io_in_key_2_0),
    .io_in_key_2_1(invkey_io_in_key_2_1),
    .io_in_key_2_2(invkey_io_in_key_2_2),
    .io_in_key_2_3(invkey_io_in_key_2_3),
    .io_in_key_3_0(invkey_io_in_key_3_0),
    .io_in_key_3_1(invkey_io_in_key_3_1),
    .io_in_key_3_2(invkey_io_in_key_3_2),
    .io_in_key_3_3(invkey_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 151:27]
  assign io_out_bits_state_0_0 = invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_1 = invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_2 = invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_3 = invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_0 = invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_1 = invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_2 = invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_3 = invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_0 = invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_1 = invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_2 = invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_3 = invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_0 = invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_1 = invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_2 = invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_3 = invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_0 = invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_1 = invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_2 = invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_3 = invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_0 = invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_1 = invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_2 = invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_3 = invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_0 = invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_1 = invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_2 = invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_3 = invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_0 = invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_1 = invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_2 = invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_3 = invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 150:18]
  assign xor__io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign sub_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign invxor_io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invmix_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invshift_io_in_state_0_0 = invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_1 = invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_2 = invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_3 = invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_0 = invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_1 = invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_2 = invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_3 = invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_0 = invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_1 = invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_2 = invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_3 = invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_0 = invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_1 = invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_2 = invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_3 = invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invsub_io_in_state_0_0 = invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_1 = invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_2 = invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_3 = invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_0 = invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_1 = invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_2 = invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_3 = invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_0 = invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_1 = invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_2 = invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_3 = invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_0 = invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_1 = invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_2 = invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_3 = invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 146:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 146:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 165:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 159:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_8(
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 237:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 240:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 241:13]
endmodule
module AES_InvGetNewKey_8(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] w4 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w5 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w6 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [31:0] w7 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] w3 = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  wire [31:0] w2 = w6 ^ w5; // @[AES_PipelinedElasticBuffer.scala 301:12]
  wire [31:0] w1 = w5 ^ w4; // @[AES_PipelinedElasticBuffer.scala 302:12]
  wire [31:0] temp = 32'h2000000 ^ sub_io_out; // @[AES_PipelinedElasticBuffer.scala 310:16]
  wire [31:0] w0 = w4 ^ temp; // @[AES_PipelinedElasticBuffer.scala 303:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 305:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 308:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w0[31:24]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_1 = w0[23:16]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_2 = w0[15:8]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_3 = w0[7:0]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_1_0 = w1[31:24]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_1 = w1[23:16]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_2 = w1[15:8]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_3 = w1[7:0]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_2_0 = w2[31:24]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_1 = w2[23:16]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_2 = w2[15:8]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_3 = w2[7:0]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_3_0 = w3[31:24]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_1 = w3[23:16]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_2 = w3[15:8]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_3 = w3[7:0]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign rot_io_in = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 309:13]
endmodule
module AES_ProcessingElement_8(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 146:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:23 AES_PipelinedElasticBuffer.scala 156:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 163:21 AES_PipelinedElasticBuffer.scala 163:21]
  AES_XOR xor_ ( // @[AES_PipelinedElasticBuffer.scala 169:19]
    .io_out_state_0_0(xor__io_out_state_0_0),
    .io_out_state_0_1(xor__io_out_state_0_1),
    .io_out_state_0_2(xor__io_out_state_0_2),
    .io_out_state_0_3(xor__io_out_state_0_3),
    .io_out_state_1_0(xor__io_out_state_1_0),
    .io_out_state_1_1(xor__io_out_state_1_1),
    .io_out_state_1_2(xor__io_out_state_1_2),
    .io_out_state_1_3(xor__io_out_state_1_3),
    .io_out_state_2_0(xor__io_out_state_2_0),
    .io_out_state_2_1(xor__io_out_state_2_1),
    .io_out_state_2_2(xor__io_out_state_2_2),
    .io_out_state_2_3(xor__io_out_state_2_3),
    .io_out_state_3_0(xor__io_out_state_3_0),
    .io_out_state_3_1(xor__io_out_state_3_1),
    .io_out_state_3_2(xor__io_out_state_3_2),
    .io_out_state_3_3(xor__io_out_state_3_3),
    .io_in_state_0_0(xor__io_in_state_0_0),
    .io_in_state_0_1(xor__io_in_state_0_1),
    .io_in_state_0_2(xor__io_in_state_0_2),
    .io_in_state_0_3(xor__io_in_state_0_3),
    .io_in_state_1_0(xor__io_in_state_1_0),
    .io_in_state_1_1(xor__io_in_state_1_1),
    .io_in_state_1_2(xor__io_in_state_1_2),
    .io_in_state_1_3(xor__io_in_state_1_3),
    .io_in_state_2_0(xor__io_in_state_2_0),
    .io_in_state_2_1(xor__io_in_state_2_1),
    .io_in_state_2_2(xor__io_in_state_2_2),
    .io_in_state_2_3(xor__io_in_state_2_3),
    .io_in_state_3_0(xor__io_in_state_3_0),
    .io_in_state_3_1(xor__io_in_state_3_1),
    .io_in_state_3_2(xor__io_in_state_3_2),
    .io_in_state_3_3(xor__io_in_state_3_3),
    .io_in_key_0_0(xor__io_in_key_0_0),
    .io_in_key_0_1(xor__io_in_key_0_1),
    .io_in_key_0_2(xor__io_in_key_0_2),
    .io_in_key_0_3(xor__io_in_key_0_3),
    .io_in_key_1_0(xor__io_in_key_1_0),
    .io_in_key_1_1(xor__io_in_key_1_1),
    .io_in_key_1_2(xor__io_in_key_1_2),
    .io_in_key_1_3(xor__io_in_key_1_3),
    .io_in_key_2_0(xor__io_in_key_2_0),
    .io_in_key_2_1(xor__io_in_key_2_1),
    .io_in_key_2_2(xor__io_in_key_2_2),
    .io_in_key_2_3(xor__io_in_key_2_3),
    .io_in_key_3_0(xor__io_in_key_3_0),
    .io_in_key_3_1(xor__io_in_key_3_1),
    .io_in_key_3_2(xor__io_in_key_3_2),
    .io_in_key_3_3(xor__io_in_key_3_3)
  );
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 174:19]
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_XOR invxor ( // @[AES_PipelinedElasticBuffer.scala 184:22]
    .io_out_state_0_0(invxor_io_out_state_0_0),
    .io_out_state_0_1(invxor_io_out_state_0_1),
    .io_out_state_0_2(invxor_io_out_state_0_2),
    .io_out_state_0_3(invxor_io_out_state_0_3),
    .io_out_state_1_0(invxor_io_out_state_1_0),
    .io_out_state_1_1(invxor_io_out_state_1_1),
    .io_out_state_1_2(invxor_io_out_state_1_2),
    .io_out_state_1_3(invxor_io_out_state_1_3),
    .io_out_state_2_0(invxor_io_out_state_2_0),
    .io_out_state_2_1(invxor_io_out_state_2_1),
    .io_out_state_2_2(invxor_io_out_state_2_2),
    .io_out_state_2_3(invxor_io_out_state_2_3),
    .io_out_state_3_0(invxor_io_out_state_3_0),
    .io_out_state_3_1(invxor_io_out_state_3_1),
    .io_out_state_3_2(invxor_io_out_state_3_2),
    .io_out_state_3_3(invxor_io_out_state_3_3),
    .io_in_state_0_0(invxor_io_in_state_0_0),
    .io_in_state_0_1(invxor_io_in_state_0_1),
    .io_in_state_0_2(invxor_io_in_state_0_2),
    .io_in_state_0_3(invxor_io_in_state_0_3),
    .io_in_state_1_0(invxor_io_in_state_1_0),
    .io_in_state_1_1(invxor_io_in_state_1_1),
    .io_in_state_1_2(invxor_io_in_state_1_2),
    .io_in_state_1_3(invxor_io_in_state_1_3),
    .io_in_state_2_0(invxor_io_in_state_2_0),
    .io_in_state_2_1(invxor_io_in_state_2_1),
    .io_in_state_2_2(invxor_io_in_state_2_2),
    .io_in_state_2_3(invxor_io_in_state_2_3),
    .io_in_state_3_0(invxor_io_in_state_3_0),
    .io_in_state_3_1(invxor_io_in_state_3_1),
    .io_in_state_3_2(invxor_io_in_state_3_2),
    .io_in_state_3_3(invxor_io_in_state_3_3),
    .io_in_key_0_0(invxor_io_in_key_0_0),
    .io_in_key_0_1(invxor_io_in_key_0_1),
    .io_in_key_0_2(invxor_io_in_key_0_2),
    .io_in_key_0_3(invxor_io_in_key_0_3),
    .io_in_key_1_0(invxor_io_in_key_1_0),
    .io_in_key_1_1(invxor_io_in_key_1_1),
    .io_in_key_1_2(invxor_io_in_key_1_2),
    .io_in_key_1_3(invxor_io_in_key_1_3),
    .io_in_key_2_0(invxor_io_in_key_2_0),
    .io_in_key_2_1(invxor_io_in_key_2_1),
    .io_in_key_2_2(invxor_io_in_key_2_2),
    .io_in_key_2_3(invxor_io_in_key_2_3),
    .io_in_key_3_0(invxor_io_in_key_3_0),
    .io_in_key_3_1(invxor_io_in_key_3_1),
    .io_in_key_3_2(invxor_io_in_key_3_2),
    .io_in_key_3_3(invxor_io_in_key_3_3)
  );
  AES_InvMixColumns invmix ( // @[AES_PipelinedElasticBuffer.scala 189:22]
    .io_out_state_0_0(invmix_io_out_state_0_0),
    .io_out_state_0_1(invmix_io_out_state_0_1),
    .io_out_state_0_2(invmix_io_out_state_0_2),
    .io_out_state_0_3(invmix_io_out_state_0_3),
    .io_out_state_1_0(invmix_io_out_state_1_0),
    .io_out_state_1_1(invmix_io_out_state_1_1),
    .io_out_state_1_2(invmix_io_out_state_1_2),
    .io_out_state_1_3(invmix_io_out_state_1_3),
    .io_out_state_2_0(invmix_io_out_state_2_0),
    .io_out_state_2_1(invmix_io_out_state_2_1),
    .io_out_state_2_2(invmix_io_out_state_2_2),
    .io_out_state_2_3(invmix_io_out_state_2_3),
    .io_out_state_3_0(invmix_io_out_state_3_0),
    .io_out_state_3_1(invmix_io_out_state_3_1),
    .io_out_state_3_2(invmix_io_out_state_3_2),
    .io_out_state_3_3(invmix_io_out_state_3_3),
    .io_in_state_0_0(invmix_io_in_state_0_0),
    .io_in_state_0_1(invmix_io_in_state_0_1),
    .io_in_state_0_2(invmix_io_in_state_0_2),
    .io_in_state_0_3(invmix_io_in_state_0_3),
    .io_in_state_1_0(invmix_io_in_state_1_0),
    .io_in_state_1_1(invmix_io_in_state_1_1),
    .io_in_state_1_2(invmix_io_in_state_1_2),
    .io_in_state_1_3(invmix_io_in_state_1_3),
    .io_in_state_2_0(invmix_io_in_state_2_0),
    .io_in_state_2_1(invmix_io_in_state_2_1),
    .io_in_state_2_2(invmix_io_in_state_2_2),
    .io_in_state_2_3(invmix_io_in_state_2_3),
    .io_in_state_3_0(invmix_io_in_state_3_0),
    .io_in_state_3_1(invmix_io_in_state_3_1),
    .io_in_state_3_2(invmix_io_in_state_3_2),
    .io_in_state_3_3(invmix_io_in_state_3_3)
  );
  AES_InvShiftRows invshift ( // @[AES_PipelinedElasticBuffer.scala 192:24]
    .io_out_state_0_0(invshift_io_out_state_0_0),
    .io_out_state_0_1(invshift_io_out_state_0_1),
    .io_out_state_0_2(invshift_io_out_state_0_2),
    .io_out_state_0_3(invshift_io_out_state_0_3),
    .io_out_state_1_0(invshift_io_out_state_1_0),
    .io_out_state_1_1(invshift_io_out_state_1_1),
    .io_out_state_1_2(invshift_io_out_state_1_2),
    .io_out_state_1_3(invshift_io_out_state_1_3),
    .io_out_state_2_0(invshift_io_out_state_2_0),
    .io_out_state_2_1(invshift_io_out_state_2_1),
    .io_out_state_2_2(invshift_io_out_state_2_2),
    .io_out_state_2_3(invshift_io_out_state_2_3),
    .io_out_state_3_0(invshift_io_out_state_3_0),
    .io_out_state_3_1(invshift_io_out_state_3_1),
    .io_out_state_3_2(invshift_io_out_state_3_2),
    .io_out_state_3_3(invshift_io_out_state_3_3),
    .io_in_state_0_0(invshift_io_in_state_0_0),
    .io_in_state_0_1(invshift_io_in_state_0_1),
    .io_in_state_0_2(invshift_io_in_state_0_2),
    .io_in_state_0_3(invshift_io_in_state_0_3),
    .io_in_state_1_0(invshift_io_in_state_1_0),
    .io_in_state_1_1(invshift_io_in_state_1_1),
    .io_in_state_1_2(invshift_io_in_state_1_2),
    .io_in_state_1_3(invshift_io_in_state_1_3),
    .io_in_state_2_0(invshift_io_in_state_2_0),
    .io_in_state_2_1(invshift_io_in_state_2_1),
    .io_in_state_2_2(invshift_io_in_state_2_2),
    .io_in_state_2_3(invshift_io_in_state_2_3),
    .io_in_state_3_0(invshift_io_in_state_3_0),
    .io_in_state_3_1(invshift_io_in_state_3_1),
    .io_in_state_3_2(invshift_io_in_state_3_2),
    .io_in_state_3_3(invshift_io_in_state_3_3)
  );
  AES_InvSubBytes invsub ( // @[AES_PipelinedElasticBuffer.scala 199:22]
    .io_out_state_0_0(invsub_io_out_state_0_0),
    .io_out_state_0_1(invsub_io_out_state_0_1),
    .io_out_state_0_2(invsub_io_out_state_0_2),
    .io_out_state_0_3(invsub_io_out_state_0_3),
    .io_out_state_1_0(invsub_io_out_state_1_0),
    .io_out_state_1_1(invsub_io_out_state_1_1),
    .io_out_state_1_2(invsub_io_out_state_1_2),
    .io_out_state_1_3(invsub_io_out_state_1_3),
    .io_out_state_2_0(invsub_io_out_state_2_0),
    .io_out_state_2_1(invsub_io_out_state_2_1),
    .io_out_state_2_2(invsub_io_out_state_2_2),
    .io_out_state_2_3(invsub_io_out_state_2_3),
    .io_out_state_3_0(invsub_io_out_state_3_0),
    .io_out_state_3_1(invsub_io_out_state_3_1),
    .io_out_state_3_2(invsub_io_out_state_3_2),
    .io_out_state_3_3(invsub_io_out_state_3_3),
    .io_in_state_0_0(invsub_io_in_state_0_0),
    .io_in_state_0_1(invsub_io_in_state_0_1),
    .io_in_state_0_2(invsub_io_in_state_0_2),
    .io_in_state_0_3(invsub_io_in_state_0_3),
    .io_in_state_1_0(invsub_io_in_state_1_0),
    .io_in_state_1_1(invsub_io_in_state_1_1),
    .io_in_state_1_2(invsub_io_in_state_1_2),
    .io_in_state_1_3(invsub_io_in_state_1_3),
    .io_in_state_2_0(invsub_io_in_state_2_0),
    .io_in_state_2_1(invsub_io_in_state_2_1),
    .io_in_state_2_2(invsub_io_in_state_2_2),
    .io_in_state_2_3(invsub_io_in_state_2_3),
    .io_in_state_3_0(invsub_io_in_state_3_0),
    .io_in_state_3_1(invsub_io_in_state_3_1),
    .io_in_state_3_2(invsub_io_in_state_3_2),
    .io_in_state_3_3(invsub_io_in_state_3_3)
  );
  AES_GetNewKey_8 key ( // @[AES_PipelinedElasticBuffer.scala 202:19]
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  AES_InvGetNewKey_8 invkey ( // @[AES_PipelinedElasticBuffer.scala 206:22]
    .io_out_key_0_0(invkey_io_out_key_0_0),
    .io_out_key_0_1(invkey_io_out_key_0_1),
    .io_out_key_0_2(invkey_io_out_key_0_2),
    .io_out_key_0_3(invkey_io_out_key_0_3),
    .io_out_key_1_0(invkey_io_out_key_1_0),
    .io_out_key_1_1(invkey_io_out_key_1_1),
    .io_out_key_1_2(invkey_io_out_key_1_2),
    .io_out_key_1_3(invkey_io_out_key_1_3),
    .io_out_key_2_0(invkey_io_out_key_2_0),
    .io_out_key_2_1(invkey_io_out_key_2_1),
    .io_out_key_2_2(invkey_io_out_key_2_2),
    .io_out_key_2_3(invkey_io_out_key_2_3),
    .io_out_key_3_0(invkey_io_out_key_3_0),
    .io_out_key_3_1(invkey_io_out_key_3_1),
    .io_out_key_3_2(invkey_io_out_key_3_2),
    .io_out_key_3_3(invkey_io_out_key_3_3),
    .io_in_key_0_0(invkey_io_in_key_0_0),
    .io_in_key_0_1(invkey_io_in_key_0_1),
    .io_in_key_0_2(invkey_io_in_key_0_2),
    .io_in_key_0_3(invkey_io_in_key_0_3),
    .io_in_key_1_0(invkey_io_in_key_1_0),
    .io_in_key_1_1(invkey_io_in_key_1_1),
    .io_in_key_1_2(invkey_io_in_key_1_2),
    .io_in_key_1_3(invkey_io_in_key_1_3),
    .io_in_key_2_0(invkey_io_in_key_2_0),
    .io_in_key_2_1(invkey_io_in_key_2_1),
    .io_in_key_2_2(invkey_io_in_key_2_2),
    .io_in_key_2_3(invkey_io_in_key_2_3),
    .io_in_key_3_0(invkey_io_in_key_3_0),
    .io_in_key_3_1(invkey_io_in_key_3_1),
    .io_in_key_3_2(invkey_io_in_key_3_2),
    .io_in_key_3_3(invkey_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 151:27]
  assign io_out_bits_state_0_0 = invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_1 = invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_2 = invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_3 = invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_0 = invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_1 = invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_2 = invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_3 = invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_0 = invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_1 = invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_2 = invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_3 = invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_0 = invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_1 = invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_2 = invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_3 = invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_0 = invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_1 = invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_2 = invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_3 = invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_0 = invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_1 = invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_2 = invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_3 = invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_0 = invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_1 = invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_2 = invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_3 = invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_0 = invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_1 = invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_2 = invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_3 = invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 150:18]
  assign xor__io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign sub_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign invxor_io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invmix_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invshift_io_in_state_0_0 = invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_1 = invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_2 = invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_3 = invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_0 = invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_1 = invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_2 = invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_3 = invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_0 = invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_1 = invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_2 = invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_3 = invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_0 = invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_1 = invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_2 = invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_3 = invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invsub_io_in_state_0_0 = invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_1 = invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_2 = invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_3 = invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_0 = invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_1 = invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_2 = invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_3 = invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_0 = invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_1 = invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_2 = invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_3 = invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_0 = invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_1 = invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_2 = invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_3 = invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 146:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 146:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 165:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 159:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_9(
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 237:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 240:19]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 237:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 240:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 241:13]
endmodule
module AES_InvGetNewKey_9(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 305:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 308:19]
  wire [31:0] w4 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w5 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w6 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [31:0] w7 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] w3 = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  wire [31:0] w2 = w6 ^ w5; // @[AES_PipelinedElasticBuffer.scala 301:12]
  wire [31:0] w1 = w5 ^ w4; // @[AES_PipelinedElasticBuffer.scala 302:12]
  wire [31:0] temp = 32'h1000000 ^ sub_io_out; // @[AES_PipelinedElasticBuffer.scala 310:16]
  wire [31:0] w0 = w4 ^ temp; // @[AES_PipelinedElasticBuffer.scala 303:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 305:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 308:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w0[31:24]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_1 = w0[23:16]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_2 = w0[15:8]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_0_3 = w0[7:0]; // @[AES_PipelinedElasticBuffer.scala 313:29]
  assign io_out_key_1_0 = w1[31:24]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_1 = w1[23:16]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_2 = w1[15:8]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_1_3 = w1[7:0]; // @[AES_PipelinedElasticBuffer.scala 314:29]
  assign io_out_key_2_0 = w2[31:24]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_1 = w2[23:16]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_2 = w2[15:8]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_2_3 = w2[7:0]; // @[AES_PipelinedElasticBuffer.scala 315:29]
  assign io_out_key_3_0 = w3[31:24]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_1 = w3[23:16]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_2 = w3[15:8]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign io_out_key_3_3 = w3[7:0]; // @[AES_PipelinedElasticBuffer.scala 316:29]
  assign rot_io_in = w7 ^ w6; // @[AES_PipelinedElasticBuffer.scala 300:12]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 309:13]
endmodule
module AES_ProcessingElement_9(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] xor__io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 169:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 174:19]
  wire [7:0] invxor_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invxor_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 184:22]
  wire [7:0] invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invmix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 189:22]
  wire [7:0] invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invshift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 192:24]
  wire [7:0] invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] invsub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 199:22]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 202:19]
  wire [7:0] invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 206:22]
  wire [7:0] invkey_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 206:22]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 145:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 146:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:23 AES_PipelinedElasticBuffer.scala 156:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 157:16 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 156:36 AES_PipelinedElasticBuffer.scala 148:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 163:21 AES_PipelinedElasticBuffer.scala 163:21]
  AES_XOR xor_ ( // @[AES_PipelinedElasticBuffer.scala 169:19]
    .io_out_state_0_0(xor__io_out_state_0_0),
    .io_out_state_0_1(xor__io_out_state_0_1),
    .io_out_state_0_2(xor__io_out_state_0_2),
    .io_out_state_0_3(xor__io_out_state_0_3),
    .io_out_state_1_0(xor__io_out_state_1_0),
    .io_out_state_1_1(xor__io_out_state_1_1),
    .io_out_state_1_2(xor__io_out_state_1_2),
    .io_out_state_1_3(xor__io_out_state_1_3),
    .io_out_state_2_0(xor__io_out_state_2_0),
    .io_out_state_2_1(xor__io_out_state_2_1),
    .io_out_state_2_2(xor__io_out_state_2_2),
    .io_out_state_2_3(xor__io_out_state_2_3),
    .io_out_state_3_0(xor__io_out_state_3_0),
    .io_out_state_3_1(xor__io_out_state_3_1),
    .io_out_state_3_2(xor__io_out_state_3_2),
    .io_out_state_3_3(xor__io_out_state_3_3),
    .io_in_state_0_0(xor__io_in_state_0_0),
    .io_in_state_0_1(xor__io_in_state_0_1),
    .io_in_state_0_2(xor__io_in_state_0_2),
    .io_in_state_0_3(xor__io_in_state_0_3),
    .io_in_state_1_0(xor__io_in_state_1_0),
    .io_in_state_1_1(xor__io_in_state_1_1),
    .io_in_state_1_2(xor__io_in_state_1_2),
    .io_in_state_1_3(xor__io_in_state_1_3),
    .io_in_state_2_0(xor__io_in_state_2_0),
    .io_in_state_2_1(xor__io_in_state_2_1),
    .io_in_state_2_2(xor__io_in_state_2_2),
    .io_in_state_2_3(xor__io_in_state_2_3),
    .io_in_state_3_0(xor__io_in_state_3_0),
    .io_in_state_3_1(xor__io_in_state_3_1),
    .io_in_state_3_2(xor__io_in_state_3_2),
    .io_in_state_3_3(xor__io_in_state_3_3),
    .io_in_key_0_0(xor__io_in_key_0_0),
    .io_in_key_0_1(xor__io_in_key_0_1),
    .io_in_key_0_2(xor__io_in_key_0_2),
    .io_in_key_0_3(xor__io_in_key_0_3),
    .io_in_key_1_0(xor__io_in_key_1_0),
    .io_in_key_1_1(xor__io_in_key_1_1),
    .io_in_key_1_2(xor__io_in_key_1_2),
    .io_in_key_1_3(xor__io_in_key_1_3),
    .io_in_key_2_0(xor__io_in_key_2_0),
    .io_in_key_2_1(xor__io_in_key_2_1),
    .io_in_key_2_2(xor__io_in_key_2_2),
    .io_in_key_2_3(xor__io_in_key_2_3),
    .io_in_key_3_0(xor__io_in_key_3_0),
    .io_in_key_3_1(xor__io_in_key_3_1),
    .io_in_key_3_2(xor__io_in_key_3_2),
    .io_in_key_3_3(xor__io_in_key_3_3)
  );
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 174:19]
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_XOR invxor ( // @[AES_PipelinedElasticBuffer.scala 184:22]
    .io_out_state_0_0(invxor_io_out_state_0_0),
    .io_out_state_0_1(invxor_io_out_state_0_1),
    .io_out_state_0_2(invxor_io_out_state_0_2),
    .io_out_state_0_3(invxor_io_out_state_0_3),
    .io_out_state_1_0(invxor_io_out_state_1_0),
    .io_out_state_1_1(invxor_io_out_state_1_1),
    .io_out_state_1_2(invxor_io_out_state_1_2),
    .io_out_state_1_3(invxor_io_out_state_1_3),
    .io_out_state_2_0(invxor_io_out_state_2_0),
    .io_out_state_2_1(invxor_io_out_state_2_1),
    .io_out_state_2_2(invxor_io_out_state_2_2),
    .io_out_state_2_3(invxor_io_out_state_2_3),
    .io_out_state_3_0(invxor_io_out_state_3_0),
    .io_out_state_3_1(invxor_io_out_state_3_1),
    .io_out_state_3_2(invxor_io_out_state_3_2),
    .io_out_state_3_3(invxor_io_out_state_3_3),
    .io_in_state_0_0(invxor_io_in_state_0_0),
    .io_in_state_0_1(invxor_io_in_state_0_1),
    .io_in_state_0_2(invxor_io_in_state_0_2),
    .io_in_state_0_3(invxor_io_in_state_0_3),
    .io_in_state_1_0(invxor_io_in_state_1_0),
    .io_in_state_1_1(invxor_io_in_state_1_1),
    .io_in_state_1_2(invxor_io_in_state_1_2),
    .io_in_state_1_3(invxor_io_in_state_1_3),
    .io_in_state_2_0(invxor_io_in_state_2_0),
    .io_in_state_2_1(invxor_io_in_state_2_1),
    .io_in_state_2_2(invxor_io_in_state_2_2),
    .io_in_state_2_3(invxor_io_in_state_2_3),
    .io_in_state_3_0(invxor_io_in_state_3_0),
    .io_in_state_3_1(invxor_io_in_state_3_1),
    .io_in_state_3_2(invxor_io_in_state_3_2),
    .io_in_state_3_3(invxor_io_in_state_3_3),
    .io_in_key_0_0(invxor_io_in_key_0_0),
    .io_in_key_0_1(invxor_io_in_key_0_1),
    .io_in_key_0_2(invxor_io_in_key_0_2),
    .io_in_key_0_3(invxor_io_in_key_0_3),
    .io_in_key_1_0(invxor_io_in_key_1_0),
    .io_in_key_1_1(invxor_io_in_key_1_1),
    .io_in_key_1_2(invxor_io_in_key_1_2),
    .io_in_key_1_3(invxor_io_in_key_1_3),
    .io_in_key_2_0(invxor_io_in_key_2_0),
    .io_in_key_2_1(invxor_io_in_key_2_1),
    .io_in_key_2_2(invxor_io_in_key_2_2),
    .io_in_key_2_3(invxor_io_in_key_2_3),
    .io_in_key_3_0(invxor_io_in_key_3_0),
    .io_in_key_3_1(invxor_io_in_key_3_1),
    .io_in_key_3_2(invxor_io_in_key_3_2),
    .io_in_key_3_3(invxor_io_in_key_3_3)
  );
  AES_InvMixColumns invmix ( // @[AES_PipelinedElasticBuffer.scala 189:22]
    .io_out_state_0_0(invmix_io_out_state_0_0),
    .io_out_state_0_1(invmix_io_out_state_0_1),
    .io_out_state_0_2(invmix_io_out_state_0_2),
    .io_out_state_0_3(invmix_io_out_state_0_3),
    .io_out_state_1_0(invmix_io_out_state_1_0),
    .io_out_state_1_1(invmix_io_out_state_1_1),
    .io_out_state_1_2(invmix_io_out_state_1_2),
    .io_out_state_1_3(invmix_io_out_state_1_3),
    .io_out_state_2_0(invmix_io_out_state_2_0),
    .io_out_state_2_1(invmix_io_out_state_2_1),
    .io_out_state_2_2(invmix_io_out_state_2_2),
    .io_out_state_2_3(invmix_io_out_state_2_3),
    .io_out_state_3_0(invmix_io_out_state_3_0),
    .io_out_state_3_1(invmix_io_out_state_3_1),
    .io_out_state_3_2(invmix_io_out_state_3_2),
    .io_out_state_3_3(invmix_io_out_state_3_3),
    .io_in_state_0_0(invmix_io_in_state_0_0),
    .io_in_state_0_1(invmix_io_in_state_0_1),
    .io_in_state_0_2(invmix_io_in_state_0_2),
    .io_in_state_0_3(invmix_io_in_state_0_3),
    .io_in_state_1_0(invmix_io_in_state_1_0),
    .io_in_state_1_1(invmix_io_in_state_1_1),
    .io_in_state_1_2(invmix_io_in_state_1_2),
    .io_in_state_1_3(invmix_io_in_state_1_3),
    .io_in_state_2_0(invmix_io_in_state_2_0),
    .io_in_state_2_1(invmix_io_in_state_2_1),
    .io_in_state_2_2(invmix_io_in_state_2_2),
    .io_in_state_2_3(invmix_io_in_state_2_3),
    .io_in_state_3_0(invmix_io_in_state_3_0),
    .io_in_state_3_1(invmix_io_in_state_3_1),
    .io_in_state_3_2(invmix_io_in_state_3_2),
    .io_in_state_3_3(invmix_io_in_state_3_3)
  );
  AES_InvShiftRows invshift ( // @[AES_PipelinedElasticBuffer.scala 192:24]
    .io_out_state_0_0(invshift_io_out_state_0_0),
    .io_out_state_0_1(invshift_io_out_state_0_1),
    .io_out_state_0_2(invshift_io_out_state_0_2),
    .io_out_state_0_3(invshift_io_out_state_0_3),
    .io_out_state_1_0(invshift_io_out_state_1_0),
    .io_out_state_1_1(invshift_io_out_state_1_1),
    .io_out_state_1_2(invshift_io_out_state_1_2),
    .io_out_state_1_3(invshift_io_out_state_1_3),
    .io_out_state_2_0(invshift_io_out_state_2_0),
    .io_out_state_2_1(invshift_io_out_state_2_1),
    .io_out_state_2_2(invshift_io_out_state_2_2),
    .io_out_state_2_3(invshift_io_out_state_2_3),
    .io_out_state_3_0(invshift_io_out_state_3_0),
    .io_out_state_3_1(invshift_io_out_state_3_1),
    .io_out_state_3_2(invshift_io_out_state_3_2),
    .io_out_state_3_3(invshift_io_out_state_3_3),
    .io_in_state_0_0(invshift_io_in_state_0_0),
    .io_in_state_0_1(invshift_io_in_state_0_1),
    .io_in_state_0_2(invshift_io_in_state_0_2),
    .io_in_state_0_3(invshift_io_in_state_0_3),
    .io_in_state_1_0(invshift_io_in_state_1_0),
    .io_in_state_1_1(invshift_io_in_state_1_1),
    .io_in_state_1_2(invshift_io_in_state_1_2),
    .io_in_state_1_3(invshift_io_in_state_1_3),
    .io_in_state_2_0(invshift_io_in_state_2_0),
    .io_in_state_2_1(invshift_io_in_state_2_1),
    .io_in_state_2_2(invshift_io_in_state_2_2),
    .io_in_state_2_3(invshift_io_in_state_2_3),
    .io_in_state_3_0(invshift_io_in_state_3_0),
    .io_in_state_3_1(invshift_io_in_state_3_1),
    .io_in_state_3_2(invshift_io_in_state_3_2),
    .io_in_state_3_3(invshift_io_in_state_3_3)
  );
  AES_InvSubBytes invsub ( // @[AES_PipelinedElasticBuffer.scala 199:22]
    .io_out_state_0_0(invsub_io_out_state_0_0),
    .io_out_state_0_1(invsub_io_out_state_0_1),
    .io_out_state_0_2(invsub_io_out_state_0_2),
    .io_out_state_0_3(invsub_io_out_state_0_3),
    .io_out_state_1_0(invsub_io_out_state_1_0),
    .io_out_state_1_1(invsub_io_out_state_1_1),
    .io_out_state_1_2(invsub_io_out_state_1_2),
    .io_out_state_1_3(invsub_io_out_state_1_3),
    .io_out_state_2_0(invsub_io_out_state_2_0),
    .io_out_state_2_1(invsub_io_out_state_2_1),
    .io_out_state_2_2(invsub_io_out_state_2_2),
    .io_out_state_2_3(invsub_io_out_state_2_3),
    .io_out_state_3_0(invsub_io_out_state_3_0),
    .io_out_state_3_1(invsub_io_out_state_3_1),
    .io_out_state_3_2(invsub_io_out_state_3_2),
    .io_out_state_3_3(invsub_io_out_state_3_3),
    .io_in_state_0_0(invsub_io_in_state_0_0),
    .io_in_state_0_1(invsub_io_in_state_0_1),
    .io_in_state_0_2(invsub_io_in_state_0_2),
    .io_in_state_0_3(invsub_io_in_state_0_3),
    .io_in_state_1_0(invsub_io_in_state_1_0),
    .io_in_state_1_1(invsub_io_in_state_1_1),
    .io_in_state_1_2(invsub_io_in_state_1_2),
    .io_in_state_1_3(invsub_io_in_state_1_3),
    .io_in_state_2_0(invsub_io_in_state_2_0),
    .io_in_state_2_1(invsub_io_in_state_2_1),
    .io_in_state_2_2(invsub_io_in_state_2_2),
    .io_in_state_2_3(invsub_io_in_state_2_3),
    .io_in_state_3_0(invsub_io_in_state_3_0),
    .io_in_state_3_1(invsub_io_in_state_3_1),
    .io_in_state_3_2(invsub_io_in_state_3_2),
    .io_in_state_3_3(invsub_io_in_state_3_3)
  );
  AES_GetNewKey_9 key ( // @[AES_PipelinedElasticBuffer.scala 202:19]
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  AES_InvGetNewKey_9 invkey ( // @[AES_PipelinedElasticBuffer.scala 206:22]
    .io_out_key_0_0(invkey_io_out_key_0_0),
    .io_out_key_0_1(invkey_io_out_key_0_1),
    .io_out_key_0_2(invkey_io_out_key_0_2),
    .io_out_key_0_3(invkey_io_out_key_0_3),
    .io_out_key_1_0(invkey_io_out_key_1_0),
    .io_out_key_1_1(invkey_io_out_key_1_1),
    .io_out_key_1_2(invkey_io_out_key_1_2),
    .io_out_key_1_3(invkey_io_out_key_1_3),
    .io_out_key_2_0(invkey_io_out_key_2_0),
    .io_out_key_2_1(invkey_io_out_key_2_1),
    .io_out_key_2_2(invkey_io_out_key_2_2),
    .io_out_key_2_3(invkey_io_out_key_2_3),
    .io_out_key_3_0(invkey_io_out_key_3_0),
    .io_out_key_3_1(invkey_io_out_key_3_1),
    .io_out_key_3_2(invkey_io_out_key_3_2),
    .io_out_key_3_3(invkey_io_out_key_3_3),
    .io_in_key_0_0(invkey_io_in_key_0_0),
    .io_in_key_0_1(invkey_io_in_key_0_1),
    .io_in_key_0_2(invkey_io_in_key_0_2),
    .io_in_key_0_3(invkey_io_in_key_0_3),
    .io_in_key_1_0(invkey_io_in_key_1_0),
    .io_in_key_1_1(invkey_io_in_key_1_1),
    .io_in_key_1_2(invkey_io_in_key_1_2),
    .io_in_key_1_3(invkey_io_in_key_1_3),
    .io_in_key_2_0(invkey_io_in_key_2_0),
    .io_in_key_2_1(invkey_io_in_key_2_1),
    .io_in_key_2_2(invkey_io_in_key_2_2),
    .io_in_key_2_3(invkey_io_in_key_2_3),
    .io_in_key_3_0(invkey_io_in_key_3_0),
    .io_in_key_3_1(invkey_io_in_key_3_1),
    .io_in_key_3_2(invkey_io_in_key_3_2),
    .io_in_key_3_3(invkey_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 151:27]
  assign io_out_bits_state_0_0 = invsub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_1 = invsub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_2 = invsub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_0_3 = invsub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_0 = invsub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_1 = invsub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_2 = invsub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_1_3 = invsub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_0 = invsub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_1 = invsub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_2 = invsub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_2_3 = invsub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_0 = invsub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_1 = invsub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_2 = invsub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_state_3_3 = invsub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_0 = invkey_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_1 = invkey_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_2 = invkey_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_0_3 = invkey_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_0 = invkey_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_1 = invkey_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_2 = invkey_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_1_3 = invkey_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_0 = invkey_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_1 = invkey_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_2 = invkey_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_2_3 = invkey_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_0 = invkey_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_1 = invkey_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_2 = invkey_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_out_bits_key_3_3 = invkey_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 152:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 150:18]
  assign xor__io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign xor__io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign sub_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign sub_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 176:19]
  assign invxor_io_in_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invxor_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invmix_io_in_state_0_0 = xor__io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_1 = xor__io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_2 = xor__io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_0_3 = xor__io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_0 = xor__io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_1 = xor__io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_2 = xor__io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_1_3 = xor__io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_0 = xor__io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_1 = xor__io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_2 = xor__io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_2_3 = xor__io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_0 = xor__io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_1 = xor__io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_2 = xor__io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invmix_io_in_state_3_3 = xor__io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 190:16]
  assign invshift_io_in_state_0_0 = invmix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_1 = invmix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_2 = invmix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_0_3 = invmix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_0 = invmix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_1 = invmix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_2 = invmix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_1_3 = invmix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_0 = invmix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_1 = invmix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_2 = invmix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_2_3 = invmix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_0 = invmix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_1 = invmix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_2 = invmix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invshift_io_in_state_3_3 = invmix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 196:20]
  assign invsub_io_in_state_0_0 = invshift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_1 = invshift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_2 = invshift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_0_3 = invshift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_0 = invshift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_1 = invshift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_2 = invshift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_1_3 = invshift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_0 = invshift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_1 = invshift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_2 = invshift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_2_3 = invshift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_0 = invshift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_1 = invshift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_2 = invshift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign invsub_io_in_state_3_3 = invshift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 200:16]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  assign invkey_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 153:9 AES_PipelinedElasticBuffer.scala 153:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 145:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 145:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 158:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 158:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 146:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 146:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 165:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 156:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 159:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 163:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 164:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 164:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_PipelinedElasticBuffer(
  input          clock,
  input          reset,
  input          io_out_ready,
  output         io_out_valid,
  output [127:0] io_out_bits_text,
  output [127:0] io_out_bits_key,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits_text,
  input  [127:0] io_in_bits_key
);
  wire  initialOperation_clock; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire  initialOperation_reset; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire  initialOperation_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire  initialOperation_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [127:0] initialOperation_io_in_bits_text; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [127:0] initialOperation_io_in_bits_key; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire  initialOperation_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire  initialOperation_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire [7:0] initialOperation_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 12:32]
  wire  finalOperation_clock; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire  finalOperation_reset; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire  finalOperation_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire  finalOperation_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [127:0] finalOperation_io_out_bits_text; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [127:0] finalOperation_io_out_bits_key; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire  finalOperation_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire  finalOperation_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire [7:0] finalOperation_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 17:30]
  wire  PEs_0_clock; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_0_reset; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_0_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_0_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_0_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_0_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_0_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_1_clock; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_1_reset; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_1_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_1_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_1_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_1_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_1_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_2_clock; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_2_reset; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_2_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_2_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_2_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_2_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_2_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_3_clock; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_3_reset; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_3_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_3_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_3_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_3_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_3_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_4_clock; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_4_reset; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_4_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_4_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_4_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_4_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_4_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_5_clock; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_5_reset; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_5_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_5_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_5_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_5_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_5_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_6_clock; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_6_reset; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_6_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_6_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_6_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_6_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_6_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_7_clock; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_7_reset; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_7_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_7_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_7_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_7_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_7_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_8_clock; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_8_reset; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_8_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_8_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_8_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_8_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_8_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_9_clock; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_9_reset; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_9_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_9_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_9_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire  PEs_9_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 23:20]
  wire [7:0] PEs_9_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 23:20]
  AES_InitialOperation initialOperation ( // @[AES_PipelinedElasticBuffer.scala 12:32]
    .clock(initialOperation_clock),
    .reset(initialOperation_reset),
    .io_in_ready(initialOperation_io_in_ready),
    .io_in_valid(initialOperation_io_in_valid),
    .io_in_bits_text(initialOperation_io_in_bits_text),
    .io_in_bits_key(initialOperation_io_in_bits_key),
    .io_out_ready(initialOperation_io_out_ready),
    .io_out_valid(initialOperation_io_out_valid),
    .io_out_bits_state_0_0(initialOperation_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(initialOperation_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(initialOperation_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(initialOperation_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(initialOperation_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(initialOperation_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(initialOperation_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(initialOperation_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(initialOperation_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(initialOperation_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(initialOperation_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(initialOperation_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(initialOperation_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(initialOperation_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(initialOperation_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(initialOperation_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(initialOperation_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(initialOperation_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(initialOperation_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(initialOperation_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(initialOperation_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(initialOperation_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(initialOperation_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(initialOperation_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(initialOperation_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(initialOperation_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(initialOperation_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(initialOperation_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(initialOperation_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(initialOperation_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(initialOperation_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(initialOperation_io_out_bits_key_3_3)
  );
  AES_FinalOperation finalOperation ( // @[AES_PipelinedElasticBuffer.scala 17:30]
    .clock(finalOperation_clock),
    .reset(finalOperation_reset),
    .io_out_ready(finalOperation_io_out_ready),
    .io_out_valid(finalOperation_io_out_valid),
    .io_out_bits_text(finalOperation_io_out_bits_text),
    .io_out_bits_key(finalOperation_io_out_bits_key),
    .io_in_ready(finalOperation_io_in_ready),
    .io_in_valid(finalOperation_io_in_valid),
    .io_in_bits_state_0_0(finalOperation_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(finalOperation_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(finalOperation_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(finalOperation_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(finalOperation_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(finalOperation_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(finalOperation_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(finalOperation_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(finalOperation_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(finalOperation_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(finalOperation_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(finalOperation_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(finalOperation_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(finalOperation_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(finalOperation_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(finalOperation_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(finalOperation_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(finalOperation_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(finalOperation_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(finalOperation_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(finalOperation_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(finalOperation_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(finalOperation_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(finalOperation_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(finalOperation_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(finalOperation_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(finalOperation_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(finalOperation_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(finalOperation_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(finalOperation_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(finalOperation_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(finalOperation_io_in_bits_key_3_3)
  );
  AES_ProcessingElement PEs_0 ( // @[AES_PipelinedElasticBuffer.scala 23:20]
    .clock(PEs_0_clock),
    .reset(PEs_0_reset),
    .io_out_ready(PEs_0_io_out_ready),
    .io_out_valid(PEs_0_io_out_valid),
    .io_out_bits_state_0_0(PEs_0_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_0_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_0_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_0_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_0_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_0_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_0_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_0_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_0_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_0_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_0_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_0_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_0_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_0_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_0_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_0_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_0_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_0_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_0_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_0_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_0_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_0_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_0_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_0_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_0_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_0_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_0_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_0_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_0_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_0_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_0_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_0_io_out_bits_key_3_3),
    .io_in_ready(PEs_0_io_in_ready),
    .io_in_valid(PEs_0_io_in_valid),
    .io_in_bits_state_0_0(PEs_0_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_0_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_0_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_0_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_0_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_0_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_0_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_0_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_0_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_0_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_0_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_0_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_0_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_0_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_0_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_0_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_0_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_0_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_0_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_0_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_0_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_0_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_0_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_0_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_0_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_0_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_0_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_0_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_0_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_0_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_0_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_0_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_1 PEs_1 ( // @[AES_PipelinedElasticBuffer.scala 23:20]
    .clock(PEs_1_clock),
    .reset(PEs_1_reset),
    .io_out_ready(PEs_1_io_out_ready),
    .io_out_valid(PEs_1_io_out_valid),
    .io_out_bits_state_0_0(PEs_1_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_1_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_1_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_1_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_1_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_1_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_1_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_1_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_1_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_1_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_1_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_1_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_1_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_1_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_1_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_1_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_1_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_1_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_1_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_1_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_1_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_1_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_1_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_1_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_1_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_1_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_1_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_1_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_1_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_1_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_1_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_1_io_out_bits_key_3_3),
    .io_in_ready(PEs_1_io_in_ready),
    .io_in_valid(PEs_1_io_in_valid),
    .io_in_bits_state_0_0(PEs_1_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_1_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_1_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_1_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_1_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_1_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_1_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_1_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_1_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_1_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_1_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_1_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_1_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_1_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_1_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_1_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_1_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_1_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_1_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_1_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_1_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_1_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_1_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_1_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_1_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_1_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_1_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_1_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_1_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_1_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_1_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_1_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_2 PEs_2 ( // @[AES_PipelinedElasticBuffer.scala 23:20]
    .clock(PEs_2_clock),
    .reset(PEs_2_reset),
    .io_out_ready(PEs_2_io_out_ready),
    .io_out_valid(PEs_2_io_out_valid),
    .io_out_bits_state_0_0(PEs_2_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_2_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_2_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_2_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_2_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_2_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_2_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_2_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_2_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_2_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_2_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_2_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_2_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_2_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_2_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_2_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_2_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_2_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_2_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_2_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_2_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_2_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_2_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_2_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_2_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_2_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_2_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_2_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_2_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_2_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_2_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_2_io_out_bits_key_3_3),
    .io_in_ready(PEs_2_io_in_ready),
    .io_in_valid(PEs_2_io_in_valid),
    .io_in_bits_state_0_0(PEs_2_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_2_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_2_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_2_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_2_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_2_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_2_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_2_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_2_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_2_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_2_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_2_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_2_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_2_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_2_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_2_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_2_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_2_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_2_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_2_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_2_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_2_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_2_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_2_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_2_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_2_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_2_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_2_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_2_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_2_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_2_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_2_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_3 PEs_3 ( // @[AES_PipelinedElasticBuffer.scala 23:20]
    .clock(PEs_3_clock),
    .reset(PEs_3_reset),
    .io_out_ready(PEs_3_io_out_ready),
    .io_out_valid(PEs_3_io_out_valid),
    .io_out_bits_state_0_0(PEs_3_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_3_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_3_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_3_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_3_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_3_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_3_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_3_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_3_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_3_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_3_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_3_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_3_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_3_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_3_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_3_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_3_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_3_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_3_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_3_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_3_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_3_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_3_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_3_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_3_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_3_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_3_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_3_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_3_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_3_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_3_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_3_io_out_bits_key_3_3),
    .io_in_ready(PEs_3_io_in_ready),
    .io_in_valid(PEs_3_io_in_valid),
    .io_in_bits_state_0_0(PEs_3_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_3_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_3_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_3_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_3_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_3_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_3_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_3_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_3_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_3_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_3_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_3_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_3_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_3_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_3_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_3_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_3_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_3_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_3_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_3_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_3_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_3_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_3_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_3_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_3_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_3_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_3_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_3_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_3_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_3_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_3_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_3_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_4 PEs_4 ( // @[AES_PipelinedElasticBuffer.scala 23:20]
    .clock(PEs_4_clock),
    .reset(PEs_4_reset),
    .io_out_ready(PEs_4_io_out_ready),
    .io_out_valid(PEs_4_io_out_valid),
    .io_out_bits_state_0_0(PEs_4_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_4_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_4_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_4_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_4_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_4_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_4_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_4_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_4_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_4_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_4_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_4_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_4_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_4_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_4_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_4_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_4_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_4_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_4_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_4_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_4_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_4_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_4_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_4_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_4_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_4_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_4_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_4_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_4_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_4_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_4_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_4_io_out_bits_key_3_3),
    .io_in_ready(PEs_4_io_in_ready),
    .io_in_valid(PEs_4_io_in_valid),
    .io_in_bits_state_0_0(PEs_4_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_4_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_4_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_4_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_4_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_4_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_4_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_4_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_4_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_4_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_4_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_4_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_4_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_4_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_4_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_4_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_4_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_4_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_4_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_4_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_4_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_4_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_4_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_4_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_4_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_4_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_4_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_4_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_4_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_4_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_4_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_4_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_5 PEs_5 ( // @[AES_PipelinedElasticBuffer.scala 23:20]
    .clock(PEs_5_clock),
    .reset(PEs_5_reset),
    .io_out_ready(PEs_5_io_out_ready),
    .io_out_valid(PEs_5_io_out_valid),
    .io_out_bits_state_0_0(PEs_5_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_5_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_5_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_5_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_5_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_5_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_5_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_5_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_5_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_5_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_5_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_5_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_5_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_5_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_5_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_5_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_5_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_5_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_5_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_5_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_5_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_5_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_5_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_5_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_5_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_5_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_5_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_5_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_5_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_5_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_5_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_5_io_out_bits_key_3_3),
    .io_in_ready(PEs_5_io_in_ready),
    .io_in_valid(PEs_5_io_in_valid),
    .io_in_bits_state_0_0(PEs_5_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_5_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_5_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_5_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_5_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_5_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_5_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_5_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_5_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_5_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_5_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_5_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_5_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_5_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_5_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_5_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_5_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_5_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_5_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_5_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_5_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_5_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_5_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_5_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_5_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_5_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_5_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_5_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_5_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_5_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_5_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_5_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_6 PEs_6 ( // @[AES_PipelinedElasticBuffer.scala 23:20]
    .clock(PEs_6_clock),
    .reset(PEs_6_reset),
    .io_out_ready(PEs_6_io_out_ready),
    .io_out_valid(PEs_6_io_out_valid),
    .io_out_bits_state_0_0(PEs_6_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_6_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_6_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_6_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_6_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_6_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_6_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_6_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_6_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_6_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_6_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_6_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_6_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_6_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_6_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_6_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_6_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_6_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_6_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_6_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_6_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_6_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_6_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_6_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_6_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_6_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_6_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_6_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_6_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_6_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_6_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_6_io_out_bits_key_3_3),
    .io_in_ready(PEs_6_io_in_ready),
    .io_in_valid(PEs_6_io_in_valid),
    .io_in_bits_state_0_0(PEs_6_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_6_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_6_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_6_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_6_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_6_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_6_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_6_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_6_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_6_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_6_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_6_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_6_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_6_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_6_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_6_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_6_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_6_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_6_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_6_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_6_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_6_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_6_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_6_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_6_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_6_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_6_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_6_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_6_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_6_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_6_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_6_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_7 PEs_7 ( // @[AES_PipelinedElasticBuffer.scala 23:20]
    .clock(PEs_7_clock),
    .reset(PEs_7_reset),
    .io_out_ready(PEs_7_io_out_ready),
    .io_out_valid(PEs_7_io_out_valid),
    .io_out_bits_state_0_0(PEs_7_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_7_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_7_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_7_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_7_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_7_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_7_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_7_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_7_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_7_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_7_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_7_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_7_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_7_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_7_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_7_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_7_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_7_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_7_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_7_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_7_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_7_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_7_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_7_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_7_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_7_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_7_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_7_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_7_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_7_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_7_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_7_io_out_bits_key_3_3),
    .io_in_ready(PEs_7_io_in_ready),
    .io_in_valid(PEs_7_io_in_valid),
    .io_in_bits_state_0_0(PEs_7_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_7_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_7_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_7_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_7_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_7_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_7_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_7_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_7_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_7_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_7_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_7_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_7_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_7_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_7_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_7_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_7_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_7_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_7_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_7_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_7_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_7_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_7_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_7_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_7_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_7_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_7_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_7_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_7_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_7_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_7_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_7_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_8 PEs_8 ( // @[AES_PipelinedElasticBuffer.scala 23:20]
    .clock(PEs_8_clock),
    .reset(PEs_8_reset),
    .io_out_ready(PEs_8_io_out_ready),
    .io_out_valid(PEs_8_io_out_valid),
    .io_out_bits_state_0_0(PEs_8_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_8_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_8_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_8_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_8_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_8_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_8_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_8_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_8_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_8_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_8_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_8_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_8_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_8_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_8_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_8_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_8_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_8_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_8_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_8_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_8_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_8_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_8_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_8_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_8_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_8_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_8_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_8_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_8_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_8_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_8_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_8_io_out_bits_key_3_3),
    .io_in_ready(PEs_8_io_in_ready),
    .io_in_valid(PEs_8_io_in_valid),
    .io_in_bits_state_0_0(PEs_8_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_8_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_8_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_8_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_8_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_8_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_8_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_8_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_8_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_8_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_8_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_8_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_8_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_8_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_8_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_8_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_8_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_8_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_8_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_8_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_8_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_8_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_8_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_8_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_8_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_8_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_8_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_8_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_8_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_8_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_8_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_8_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_9 PEs_9 ( // @[AES_PipelinedElasticBuffer.scala 23:20]
    .clock(PEs_9_clock),
    .reset(PEs_9_reset),
    .io_out_ready(PEs_9_io_out_ready),
    .io_out_valid(PEs_9_io_out_valid),
    .io_out_bits_state_0_0(PEs_9_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_9_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_9_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_9_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_9_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_9_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_9_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_9_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_9_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_9_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_9_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_9_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_9_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_9_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_9_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_9_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_9_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_9_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_9_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_9_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_9_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_9_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_9_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_9_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_9_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_9_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_9_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_9_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_9_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_9_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_9_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_9_io_out_bits_key_3_3),
    .io_in_ready(PEs_9_io_in_ready),
    .io_in_valid(PEs_9_io_in_valid),
    .io_in_bits_state_0_0(PEs_9_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_9_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_9_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_9_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_9_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_9_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_9_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_9_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_9_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_9_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_9_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_9_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_9_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_9_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_9_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_9_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_9_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_9_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_9_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_9_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_9_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_9_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_9_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_9_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_9_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_9_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_9_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_9_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_9_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_9_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_9_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_9_io_in_bits_key_3_3)
  );
  assign io_out_valid = finalOperation_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 19:16]
  assign io_out_bits_text = finalOperation_io_out_bits_text; // @[AES_PipelinedElasticBuffer.scala 18:15]
  assign io_out_bits_key = finalOperation_io_out_bits_key; // @[AES_PipelinedElasticBuffer.scala 18:15]
  assign io_in_ready = initialOperation_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 15:15]
  assign initialOperation_clock = clock;
  assign initialOperation_reset = reset;
  assign initialOperation_io_in_valid = io_in_valid; // @[AES_PipelinedElasticBuffer.scala 13:32]
  assign initialOperation_io_in_bits_text = io_in_bits_text; // @[AES_PipelinedElasticBuffer.scala 14:31]
  assign initialOperation_io_in_bits_key = io_in_bits_key; // @[AES_PipelinedElasticBuffer.scala 14:31]
  assign initialOperation_io_out_ready = PEs_0_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 32:37]
  assign finalOperation_clock = clock;
  assign finalOperation_reset = reset;
  assign finalOperation_io_out_ready = io_out_ready; // @[AES_PipelinedElasticBuffer.scala 20:31]
  assign finalOperation_io_in_valid = PEs_9_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 38:34]
  assign finalOperation_io_in_bits_state_0_0 = PEs_9_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_0_1 = PEs_9_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_0_2 = PEs_9_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_0_3 = PEs_9_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_1_0 = PEs_9_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_1_1 = PEs_9_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_1_2 = PEs_9_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_1_3 = PEs_9_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_2_0 = PEs_9_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_2_1 = PEs_9_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_2_2 = PEs_9_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_2_3 = PEs_9_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_3_0 = PEs_9_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_3_1 = PEs_9_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_3_2 = PEs_9_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_state_3_3 = PEs_9_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 39:39]
  assign finalOperation_io_in_bits_key_0_0 = PEs_9_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_0_1 = PEs_9_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_0_2 = PEs_9_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_0_3 = PEs_9_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_1_0 = PEs_9_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_1_1 = PEs_9_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_1_2 = PEs_9_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_1_3 = PEs_9_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_2_0 = PEs_9_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_2_1 = PEs_9_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_2_2 = PEs_9_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_2_3 = PEs_9_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_3_0 = PEs_9_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_3_1 = PEs_9_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_3_2 = PEs_9_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign finalOperation_io_in_bits_key_3_3 = PEs_9_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 40:37]
  assign PEs_0_clock = clock;
  assign PEs_0_reset = reset;
  assign PEs_0_io_out_ready = PEs_1_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 36:27]
  assign PEs_0_io_in_valid = initialOperation_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 30:26]
  assign PEs_0_io_in_bits_state_0_0 = initialOperation_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_0_1 = initialOperation_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_0_2 = initialOperation_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_0_3 = initialOperation_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_1_0 = initialOperation_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_1_1 = initialOperation_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_1_2 = initialOperation_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_1_3 = initialOperation_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_2_0 = initialOperation_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_2_1 = initialOperation_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_2_2 = initialOperation_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_2_3 = initialOperation_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_3_0 = initialOperation_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_3_1 = initialOperation_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_3_2 = initialOperation_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_state_3_3 = initialOperation_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_0_0 = initialOperation_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_0_1 = initialOperation_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_0_2 = initialOperation_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_0_3 = initialOperation_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_1_0 = initialOperation_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_1_1 = initialOperation_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_1_2 = initialOperation_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_1_3 = initialOperation_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_2_0 = initialOperation_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_2_1 = initialOperation_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_2_2 = initialOperation_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_2_3 = initialOperation_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_3_0 = initialOperation_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_3_1 = initialOperation_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_3_2 = initialOperation_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_0_io_in_bits_key_3_3 = initialOperation_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 31:25]
  assign PEs_1_clock = clock;
  assign PEs_1_reset = reset;
  assign PEs_1_io_out_ready = PEs_2_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 45:27]
  assign PEs_1_io_in_valid = PEs_0_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 34:28]
  assign PEs_1_io_in_bits_state_0_0 = PEs_0_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_0_1 = PEs_0_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_0_2 = PEs_0_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_0_3 = PEs_0_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_1_0 = PEs_0_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_1_1 = PEs_0_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_1_2 = PEs_0_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_1_3 = PEs_0_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_2_0 = PEs_0_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_2_1 = PEs_0_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_2_2 = PEs_0_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_2_3 = PEs_0_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_3_0 = PEs_0_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_3_1 = PEs_0_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_3_2 = PEs_0_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_state_3_3 = PEs_0_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_0_0 = PEs_0_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_0_1 = PEs_0_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_0_2 = PEs_0_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_0_3 = PEs_0_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_1_0 = PEs_0_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_1_1 = PEs_0_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_1_2 = PEs_0_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_1_3 = PEs_0_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_2_0 = PEs_0_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_2_1 = PEs_0_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_2_2 = PEs_0_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_2_3 = PEs_0_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_3_0 = PEs_0_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_3_1 = PEs_0_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_3_2 = PEs_0_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_1_io_in_bits_key_3_3 = PEs_0_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 35:27]
  assign PEs_2_clock = clock;
  assign PEs_2_reset = reset;
  assign PEs_2_io_out_ready = PEs_3_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 45:27]
  assign PEs_2_io_in_valid = PEs_1_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 43:28]
  assign PEs_2_io_in_bits_state_0_0 = PEs_1_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_0_1 = PEs_1_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_0_2 = PEs_1_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_0_3 = PEs_1_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_1_0 = PEs_1_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_1_1 = PEs_1_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_1_2 = PEs_1_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_1_3 = PEs_1_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_2_0 = PEs_1_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_2_1 = PEs_1_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_2_2 = PEs_1_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_2_3 = PEs_1_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_3_0 = PEs_1_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_3_1 = PEs_1_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_3_2 = PEs_1_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_state_3_3 = PEs_1_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_0_0 = PEs_1_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_0_1 = PEs_1_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_0_2 = PEs_1_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_0_3 = PEs_1_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_1_0 = PEs_1_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_1_1 = PEs_1_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_1_2 = PEs_1_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_1_3 = PEs_1_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_2_0 = PEs_1_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_2_1 = PEs_1_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_2_2 = PEs_1_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_2_3 = PEs_1_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_3_0 = PEs_1_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_3_1 = PEs_1_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_3_2 = PEs_1_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_2_io_in_bits_key_3_3 = PEs_1_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_clock = clock;
  assign PEs_3_reset = reset;
  assign PEs_3_io_out_ready = PEs_4_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 45:27]
  assign PEs_3_io_in_valid = PEs_2_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 43:28]
  assign PEs_3_io_in_bits_state_0_0 = PEs_2_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_0_1 = PEs_2_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_0_2 = PEs_2_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_0_3 = PEs_2_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_1_0 = PEs_2_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_1_1 = PEs_2_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_1_2 = PEs_2_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_1_3 = PEs_2_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_2_0 = PEs_2_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_2_1 = PEs_2_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_2_2 = PEs_2_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_2_3 = PEs_2_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_3_0 = PEs_2_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_3_1 = PEs_2_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_3_2 = PEs_2_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_state_3_3 = PEs_2_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_0_0 = PEs_2_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_0_1 = PEs_2_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_0_2 = PEs_2_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_0_3 = PEs_2_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_1_0 = PEs_2_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_1_1 = PEs_2_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_1_2 = PEs_2_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_1_3 = PEs_2_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_2_0 = PEs_2_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_2_1 = PEs_2_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_2_2 = PEs_2_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_2_3 = PEs_2_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_3_0 = PEs_2_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_3_1 = PEs_2_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_3_2 = PEs_2_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_3_io_in_bits_key_3_3 = PEs_2_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_clock = clock;
  assign PEs_4_reset = reset;
  assign PEs_4_io_out_ready = PEs_5_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 45:27]
  assign PEs_4_io_in_valid = PEs_3_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 43:28]
  assign PEs_4_io_in_bits_state_0_0 = PEs_3_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_0_1 = PEs_3_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_0_2 = PEs_3_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_0_3 = PEs_3_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_1_0 = PEs_3_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_1_1 = PEs_3_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_1_2 = PEs_3_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_1_3 = PEs_3_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_2_0 = PEs_3_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_2_1 = PEs_3_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_2_2 = PEs_3_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_2_3 = PEs_3_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_3_0 = PEs_3_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_3_1 = PEs_3_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_3_2 = PEs_3_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_state_3_3 = PEs_3_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_0_0 = PEs_3_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_0_1 = PEs_3_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_0_2 = PEs_3_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_0_3 = PEs_3_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_1_0 = PEs_3_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_1_1 = PEs_3_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_1_2 = PEs_3_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_1_3 = PEs_3_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_2_0 = PEs_3_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_2_1 = PEs_3_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_2_2 = PEs_3_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_2_3 = PEs_3_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_3_0 = PEs_3_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_3_1 = PEs_3_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_3_2 = PEs_3_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_4_io_in_bits_key_3_3 = PEs_3_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_clock = clock;
  assign PEs_5_reset = reset;
  assign PEs_5_io_out_ready = PEs_6_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 45:27]
  assign PEs_5_io_in_valid = PEs_4_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 43:28]
  assign PEs_5_io_in_bits_state_0_0 = PEs_4_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_0_1 = PEs_4_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_0_2 = PEs_4_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_0_3 = PEs_4_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_1_0 = PEs_4_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_1_1 = PEs_4_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_1_2 = PEs_4_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_1_3 = PEs_4_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_2_0 = PEs_4_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_2_1 = PEs_4_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_2_2 = PEs_4_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_2_3 = PEs_4_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_3_0 = PEs_4_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_3_1 = PEs_4_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_3_2 = PEs_4_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_state_3_3 = PEs_4_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_0_0 = PEs_4_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_0_1 = PEs_4_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_0_2 = PEs_4_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_0_3 = PEs_4_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_1_0 = PEs_4_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_1_1 = PEs_4_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_1_2 = PEs_4_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_1_3 = PEs_4_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_2_0 = PEs_4_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_2_1 = PEs_4_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_2_2 = PEs_4_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_2_3 = PEs_4_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_3_0 = PEs_4_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_3_1 = PEs_4_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_3_2 = PEs_4_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_5_io_in_bits_key_3_3 = PEs_4_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_clock = clock;
  assign PEs_6_reset = reset;
  assign PEs_6_io_out_ready = PEs_7_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 45:27]
  assign PEs_6_io_in_valid = PEs_5_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 43:28]
  assign PEs_6_io_in_bits_state_0_0 = PEs_5_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_0_1 = PEs_5_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_0_2 = PEs_5_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_0_3 = PEs_5_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_1_0 = PEs_5_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_1_1 = PEs_5_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_1_2 = PEs_5_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_1_3 = PEs_5_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_2_0 = PEs_5_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_2_1 = PEs_5_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_2_2 = PEs_5_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_2_3 = PEs_5_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_3_0 = PEs_5_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_3_1 = PEs_5_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_3_2 = PEs_5_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_state_3_3 = PEs_5_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_0_0 = PEs_5_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_0_1 = PEs_5_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_0_2 = PEs_5_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_0_3 = PEs_5_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_1_0 = PEs_5_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_1_1 = PEs_5_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_1_2 = PEs_5_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_1_3 = PEs_5_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_2_0 = PEs_5_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_2_1 = PEs_5_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_2_2 = PEs_5_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_2_3 = PEs_5_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_3_0 = PEs_5_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_3_1 = PEs_5_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_3_2 = PEs_5_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_6_io_in_bits_key_3_3 = PEs_5_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_clock = clock;
  assign PEs_7_reset = reset;
  assign PEs_7_io_out_ready = PEs_8_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 45:27]
  assign PEs_7_io_in_valid = PEs_6_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 43:28]
  assign PEs_7_io_in_bits_state_0_0 = PEs_6_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_0_1 = PEs_6_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_0_2 = PEs_6_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_0_3 = PEs_6_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_1_0 = PEs_6_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_1_1 = PEs_6_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_1_2 = PEs_6_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_1_3 = PEs_6_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_2_0 = PEs_6_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_2_1 = PEs_6_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_2_2 = PEs_6_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_2_3 = PEs_6_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_3_0 = PEs_6_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_3_1 = PEs_6_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_3_2 = PEs_6_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_state_3_3 = PEs_6_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_0_0 = PEs_6_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_0_1 = PEs_6_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_0_2 = PEs_6_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_0_3 = PEs_6_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_1_0 = PEs_6_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_1_1 = PEs_6_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_1_2 = PEs_6_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_1_3 = PEs_6_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_2_0 = PEs_6_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_2_1 = PEs_6_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_2_2 = PEs_6_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_2_3 = PEs_6_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_3_0 = PEs_6_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_3_1 = PEs_6_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_3_2 = PEs_6_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_7_io_in_bits_key_3_3 = PEs_6_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_clock = clock;
  assign PEs_8_reset = reset;
  assign PEs_8_io_out_ready = PEs_9_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 45:27]
  assign PEs_8_io_in_valid = PEs_7_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 43:28]
  assign PEs_8_io_in_bits_state_0_0 = PEs_7_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_0_1 = PEs_7_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_0_2 = PEs_7_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_0_3 = PEs_7_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_1_0 = PEs_7_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_1_1 = PEs_7_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_1_2 = PEs_7_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_1_3 = PEs_7_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_2_0 = PEs_7_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_2_1 = PEs_7_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_2_2 = PEs_7_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_2_3 = PEs_7_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_3_0 = PEs_7_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_3_1 = PEs_7_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_3_2 = PEs_7_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_state_3_3 = PEs_7_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_0_0 = PEs_7_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_0_1 = PEs_7_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_0_2 = PEs_7_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_0_3 = PEs_7_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_1_0 = PEs_7_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_1_1 = PEs_7_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_1_2 = PEs_7_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_1_3 = PEs_7_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_2_0 = PEs_7_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_2_1 = PEs_7_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_2_2 = PEs_7_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_2_3 = PEs_7_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_3_0 = PEs_7_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_3_1 = PEs_7_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_3_2 = PEs_7_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_8_io_in_bits_key_3_3 = PEs_7_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_clock = clock;
  assign PEs_9_reset = reset;
  assign PEs_9_io_out_ready = finalOperation_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 41:27]
  assign PEs_9_io_in_valid = PEs_8_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 43:28]
  assign PEs_9_io_in_bits_state_0_0 = PEs_8_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_0_1 = PEs_8_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_0_2 = PEs_8_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_0_3 = PEs_8_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_1_0 = PEs_8_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_1_1 = PEs_8_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_1_2 = PEs_8_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_1_3 = PEs_8_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_2_0 = PEs_8_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_2_1 = PEs_8_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_2_2 = PEs_8_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_2_3 = PEs_8_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_3_0 = PEs_8_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_3_1 = PEs_8_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_3_2 = PEs_8_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_state_3_3 = PEs_8_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_0_0 = PEs_8_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_0_1 = PEs_8_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_0_2 = PEs_8_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_0_3 = PEs_8_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_1_0 = PEs_8_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_1_1 = PEs_8_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_1_2 = PEs_8_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_1_3 = PEs_8_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_2_0 = PEs_8_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_2_1 = PEs_8_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_2_2 = PEs_8_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_2_3 = PEs_8_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_3_0 = PEs_8_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_3_1 = PEs_8_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_3_2 = PEs_8_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 44:27]
  assign PEs_9_io_in_bits_key_3_3 = PEs_8_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 44:27]
endmodule
