module IP(
  input  [63:0] io_text,
  output [31:0] io_L,
  output [31:0] io_R
);
  wire [63:0] _T_3 = {{32'd0}, io_text[63:32]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_5 = {io_text[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_7 = _T_5 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_8 = _T_3 | _T_7; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_0 = {{16'd0}, _T_8[63:16]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_13 = _GEN_0 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_15 = {_T_8[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_17 = _T_15 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_18 = _T_13 | _T_17; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_1 = {{8'd0}, _T_18[63:8]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_23 = _GEN_1 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_25 = {_T_18[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_27 = _T_25 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  wire [63:0] _T_28 = _T_23 | _T_27; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_2 = {{4'd0}, _T_28[63:4]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_33 = _GEN_2 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  wire [63:0] _T_35 = {_T_28[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_37 = _T_35 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  wire [63:0] _T_38 = _T_33 | _T_37; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_3 = {{2'd0}, _T_38[63:2]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_43 = _GEN_3 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  wire [63:0] _T_45 = {_T_38[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_47 = _T_45 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  wire [63:0] _T_48 = _T_43 | _T_47; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_4 = {{1'd0}, _T_48[63:1]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_53 = _GEN_4 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  wire [63:0] _T_55 = {_T_48[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_57 = _T_55 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  wire [63:0] reversed = _T_53 | _T_57; // @[Bitwise.scala 103:39]
  wire  hi_hi_hi_hi_hi = reversed[57]; // @[DES_FSM.scala 147:23]
  wire  hi_hi_hi_hi_lo = reversed[49]; // @[DES_FSM.scala 147:36]
  wire  hi_hi_hi_lo_hi = reversed[41]; // @[DES_FSM.scala 147:49]
  wire  hi_hi_hi_lo_lo = reversed[33]; // @[DES_FSM.scala 147:62]
  wire  hi_hi_lo_hi_hi = reversed[25]; // @[DES_FSM.scala 147:75]
  wire  hi_hi_lo_hi_lo = reversed[17]; // @[DES_FSM.scala 147:88]
  wire  hi_hi_lo_lo_hi = reversed[9]; // @[DES_FSM.scala 147:101]
  wire  hi_hi_lo_lo_lo = reversed[1]; // @[DES_FSM.scala 147:113]
  wire  hi_lo_hi_hi_hi = reversed[59]; // @[DES_FSM.scala 148:13]
  wire  hi_lo_hi_hi_lo = reversed[51]; // @[DES_FSM.scala 148:26]
  wire  hi_lo_hi_lo_hi = reversed[43]; // @[DES_FSM.scala 148:39]
  wire  hi_lo_hi_lo_lo = reversed[35]; // @[DES_FSM.scala 148:52]
  wire  hi_lo_lo_hi_hi = reversed[27]; // @[DES_FSM.scala 148:65]
  wire  hi_lo_lo_hi_lo = reversed[19]; // @[DES_FSM.scala 148:78]
  wire  hi_lo_lo_lo_hi = reversed[11]; // @[DES_FSM.scala 148:91]
  wire  hi_lo_lo_lo_lo = reversed[3]; // @[DES_FSM.scala 148:104]
  wire  lo_hi_hi_hi_hi = reversed[61]; // @[DES_FSM.scala 149:13]
  wire  lo_hi_hi_hi_lo = reversed[53]; // @[DES_FSM.scala 149:26]
  wire  lo_hi_hi_lo_hi = reversed[45]; // @[DES_FSM.scala 149:39]
  wire  lo_hi_hi_lo_lo = reversed[37]; // @[DES_FSM.scala 149:52]
  wire  lo_hi_lo_hi_hi = reversed[29]; // @[DES_FSM.scala 149:65]
  wire  lo_hi_lo_hi_lo = reversed[21]; // @[DES_FSM.scala 149:78]
  wire  lo_hi_lo_lo_hi = reversed[13]; // @[DES_FSM.scala 149:91]
  wire  lo_hi_lo_lo_lo = reversed[5]; // @[DES_FSM.scala 149:104]
  wire  lo_lo_hi_hi_hi = reversed[63]; // @[DES_FSM.scala 150:13]
  wire  lo_lo_hi_hi_lo = reversed[55]; // @[DES_FSM.scala 150:26]
  wire  lo_lo_hi_lo_hi = reversed[47]; // @[DES_FSM.scala 150:39]
  wire  lo_lo_hi_lo_lo = reversed[39]; // @[DES_FSM.scala 150:52]
  wire  lo_lo_lo_hi_hi = reversed[31]; // @[DES_FSM.scala 150:65]
  wire  lo_lo_lo_hi_lo = reversed[23]; // @[DES_FSM.scala 150:78]
  wire  lo_lo_lo_lo_hi = reversed[15]; // @[DES_FSM.scala 150:91]
  wire  lo_lo_lo_lo_lo = reversed[7]; // @[DES_FSM.scala 150:104]
  wire [7:0] lo_lo = {lo_lo_hi_hi_hi,lo_lo_hi_hi_lo,lo_lo_hi_lo_hi,lo_lo_hi_lo_lo,lo_lo_lo_hi_hi,lo_lo_lo_hi_lo,
    lo_lo_lo_lo_hi,lo_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [15:0] lo = {lo_hi_hi_hi_hi,lo_hi_hi_hi_lo,lo_hi_hi_lo_hi,lo_hi_hi_lo_lo,lo_hi_lo_hi_hi,lo_hi_lo_hi_lo,
    lo_hi_lo_lo_hi,lo_hi_lo_lo_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo = {hi_lo_hi_hi_hi,hi_lo_hi_hi_lo,hi_lo_hi_lo_hi,hi_lo_hi_lo_lo,hi_lo_lo_hi_hi,hi_lo_lo_hi_lo,
    hi_lo_lo_lo_hi,hi_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [15:0] hi = {hi_hi_hi_hi_hi,hi_hi_hi_hi_lo,hi_hi_hi_lo_hi,hi_hi_hi_lo_lo,hi_hi_lo_hi_hi,hi_hi_lo_hi_lo,
    hi_hi_lo_lo_hi,hi_hi_lo_lo_lo,hi_lo}; // @[Cat.scala 30:58]
  wire  hi_hi_hi_hi_hi_1 = reversed[56]; // @[DES_FSM.scala 152:23]
  wire  hi_hi_hi_hi_lo_1 = reversed[48]; // @[DES_FSM.scala 152:36]
  wire  hi_hi_hi_lo_hi_1 = reversed[40]; // @[DES_FSM.scala 152:49]
  wire  hi_hi_hi_lo_lo_1 = reversed[32]; // @[DES_FSM.scala 152:62]
  wire  hi_hi_lo_hi_hi_1 = reversed[24]; // @[DES_FSM.scala 152:75]
  wire  hi_hi_lo_hi_lo_1 = reversed[16]; // @[DES_FSM.scala 152:88]
  wire  hi_hi_lo_lo_hi_1 = reversed[8]; // @[DES_FSM.scala 152:101]
  wire  hi_hi_lo_lo_lo_1 = reversed[0]; // @[DES_FSM.scala 152:113]
  wire  hi_lo_hi_hi_hi_1 = reversed[58]; // @[DES_FSM.scala 153:13]
  wire  hi_lo_hi_hi_lo_1 = reversed[50]; // @[DES_FSM.scala 153:26]
  wire  hi_lo_hi_lo_hi_1 = reversed[42]; // @[DES_FSM.scala 153:39]
  wire  hi_lo_hi_lo_lo_1 = reversed[34]; // @[DES_FSM.scala 153:52]
  wire  hi_lo_lo_hi_hi_1 = reversed[26]; // @[DES_FSM.scala 153:65]
  wire  hi_lo_lo_hi_lo_1 = reversed[18]; // @[DES_FSM.scala 153:78]
  wire  hi_lo_lo_lo_hi_1 = reversed[10]; // @[DES_FSM.scala 153:91]
  wire  hi_lo_lo_lo_lo_1 = reversed[2]; // @[DES_FSM.scala 153:104]
  wire  lo_hi_hi_hi_hi_1 = reversed[60]; // @[DES_FSM.scala 154:13]
  wire  lo_hi_hi_hi_lo_1 = reversed[52]; // @[DES_FSM.scala 154:26]
  wire  lo_hi_hi_lo_hi_1 = reversed[44]; // @[DES_FSM.scala 154:39]
  wire  lo_hi_hi_lo_lo_1 = reversed[36]; // @[DES_FSM.scala 154:52]
  wire  lo_hi_lo_hi_hi_1 = reversed[28]; // @[DES_FSM.scala 154:65]
  wire  lo_hi_lo_hi_lo_1 = reversed[20]; // @[DES_FSM.scala 154:78]
  wire  lo_hi_lo_lo_hi_1 = reversed[12]; // @[DES_FSM.scala 154:91]
  wire  lo_hi_lo_lo_lo_1 = reversed[4]; // @[DES_FSM.scala 154:104]
  wire  lo_lo_hi_hi_hi_1 = reversed[62]; // @[DES_FSM.scala 155:13]
  wire  lo_lo_hi_hi_lo_1 = reversed[54]; // @[DES_FSM.scala 155:26]
  wire  lo_lo_hi_lo_hi_1 = reversed[46]; // @[DES_FSM.scala 155:39]
  wire  lo_lo_hi_lo_lo_1 = reversed[38]; // @[DES_FSM.scala 155:52]
  wire  lo_lo_lo_hi_hi_1 = reversed[30]; // @[DES_FSM.scala 155:65]
  wire  lo_lo_lo_hi_lo_1 = reversed[22]; // @[DES_FSM.scala 155:78]
  wire  lo_lo_lo_lo_hi_1 = reversed[14]; // @[DES_FSM.scala 155:91]
  wire  lo_lo_lo_lo_lo_1 = reversed[6]; // @[DES_FSM.scala 155:104]
  wire [7:0] lo_lo_1 = {lo_lo_hi_hi_hi_1,lo_lo_hi_hi_lo_1,lo_lo_hi_lo_hi_1,lo_lo_hi_lo_lo_1,lo_lo_lo_hi_hi_1,
    lo_lo_lo_hi_lo_1,lo_lo_lo_lo_hi_1,lo_lo_lo_lo_lo_1}; // @[Cat.scala 30:58]
  wire [15:0] lo_1 = {lo_hi_hi_hi_hi_1,lo_hi_hi_hi_lo_1,lo_hi_hi_lo_hi_1,lo_hi_hi_lo_lo_1,lo_hi_lo_hi_hi_1,
    lo_hi_lo_hi_lo_1,lo_hi_lo_lo_hi_1,lo_hi_lo_lo_lo_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo_1 = {hi_lo_hi_hi_hi_1,hi_lo_hi_hi_lo_1,hi_lo_hi_lo_hi_1,hi_lo_hi_lo_lo_1,hi_lo_lo_hi_hi_1,
    hi_lo_lo_hi_lo_1,hi_lo_lo_lo_hi_1,hi_lo_lo_lo_lo_1}; // @[Cat.scala 30:58]
  wire [15:0] hi_1 = {hi_hi_hi_hi_hi_1,hi_hi_hi_hi_lo_1,hi_hi_hi_lo_hi_1,hi_hi_hi_lo_lo_1,hi_hi_lo_hi_hi_1,
    hi_hi_lo_hi_lo_1,hi_hi_lo_lo_hi_1,hi_hi_lo_lo_lo_1,hi_lo_1}; // @[Cat.scala 30:58]
  assign io_L = {hi,lo}; // @[Cat.scala 30:58]
  assign io_R = {hi_1,lo_1}; // @[Cat.scala 30:58]
endmodule
module PC_1(
  input  [63:0] io_key,
  output [27:0] io_C,
  output [27:0] io_D
);
  wire [63:0] _T_3 = {{32'd0}, io_key[63:32]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_5 = {io_key[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_7 = _T_5 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_8 = _T_3 | _T_7; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_0 = {{16'd0}, _T_8[63:16]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_13 = _GEN_0 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_15 = {_T_8[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_17 = _T_15 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_18 = _T_13 | _T_17; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_1 = {{8'd0}, _T_18[63:8]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_23 = _GEN_1 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_25 = {_T_18[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_27 = _T_25 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  wire [63:0] _T_28 = _T_23 | _T_27; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_2 = {{4'd0}, _T_28[63:4]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_33 = _GEN_2 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  wire [63:0] _T_35 = {_T_28[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_37 = _T_35 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  wire [63:0] _T_38 = _T_33 | _T_37; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_3 = {{2'd0}, _T_38[63:2]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_43 = _GEN_3 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  wire [63:0] _T_45 = {_T_38[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_47 = _T_45 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  wire [63:0] _T_48 = _T_43 | _T_47; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_4 = {{1'd0}, _T_48[63:1]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_53 = _GEN_4 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  wire [63:0] _T_55 = {_T_48[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_57 = _T_55 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  wire [63:0] reversed = _T_53 | _T_57; // @[Bitwise.scala 103:39]
  wire  hi_hi_hi_hi_hi = reversed[56]; // @[DES_FSM.scala 168:23]
  wire  hi_hi_hi_hi_lo = reversed[48]; // @[DES_FSM.scala 168:36]
  wire  hi_hi_hi_lo_hi = reversed[40]; // @[DES_FSM.scala 168:49]
  wire  hi_hi_hi_lo_lo = reversed[32]; // @[DES_FSM.scala 168:62]
  wire  hi_hi_lo_hi_hi = reversed[24]; // @[DES_FSM.scala 168:75]
  wire  hi_hi_lo_hi_lo = reversed[16]; // @[DES_FSM.scala 168:88]
  wire  hi_hi_lo_lo = reversed[8]; // @[DES_FSM.scala 168:101]
  wire  hi_lo_hi_hi_hi = reversed[0]; // @[DES_FSM.scala 169:13]
  wire  hi_lo_hi_hi_lo = reversed[57]; // @[DES_FSM.scala 169:25]
  wire  hi_lo_hi_lo_hi = reversed[49]; // @[DES_FSM.scala 169:38]
  wire  hi_lo_hi_lo_lo = reversed[41]; // @[DES_FSM.scala 169:51]
  wire  hi_lo_lo_hi_hi = reversed[33]; // @[DES_FSM.scala 169:64]
  wire  hi_lo_lo_hi_lo = reversed[25]; // @[DES_FSM.scala 169:77]
  wire  hi_lo_lo_lo = reversed[17]; // @[DES_FSM.scala 169:90]
  wire  lo_hi_hi_hi_hi = reversed[9]; // @[DES_FSM.scala 170:13]
  wire  lo_hi_hi_hi_lo = reversed[1]; // @[DES_FSM.scala 170:25]
  wire  lo_hi_hi_lo_hi = reversed[58]; // @[DES_FSM.scala 170:37]
  wire  lo_hi_hi_lo_lo = reversed[50]; // @[DES_FSM.scala 170:50]
  wire  lo_hi_lo_hi_hi = reversed[42]; // @[DES_FSM.scala 170:63]
  wire  lo_hi_lo_hi_lo = reversed[34]; // @[DES_FSM.scala 170:76]
  wire  lo_hi_lo_lo = reversed[26]; // @[DES_FSM.scala 170:89]
  wire  lo_lo_hi_hi_hi = reversed[18]; // @[DES_FSM.scala 171:13]
  wire  lo_lo_hi_hi_lo = reversed[10]; // @[DES_FSM.scala 171:26]
  wire  lo_lo_hi_lo_hi = reversed[2]; // @[DES_FSM.scala 171:39]
  wire  lo_lo_hi_lo_lo = reversed[59]; // @[DES_FSM.scala 171:51]
  wire  lo_lo_lo_hi_hi = reversed[51]; // @[DES_FSM.scala 171:64]
  wire  lo_lo_lo_hi_lo = reversed[43]; // @[DES_FSM.scala 171:77]
  wire  lo_lo_lo_lo = reversed[35]; // @[DES_FSM.scala 171:90]
  wire [6:0] lo_lo = {lo_lo_hi_hi_hi,lo_lo_hi_hi_lo,lo_lo_hi_lo_hi,lo_lo_hi_lo_lo,lo_lo_lo_hi_hi,lo_lo_lo_hi_lo,
    lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [13:0] lo = {lo_hi_hi_hi_hi,lo_hi_hi_hi_lo,lo_hi_hi_lo_hi,lo_hi_hi_lo_lo,lo_hi_lo_hi_hi,lo_hi_lo_hi_lo,
    lo_hi_lo_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [6:0] hi_lo = {hi_lo_hi_hi_hi,hi_lo_hi_hi_lo,hi_lo_hi_lo_hi,hi_lo_hi_lo_lo,hi_lo_lo_hi_hi,hi_lo_lo_hi_lo,
    hi_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [13:0] hi = {hi_hi_hi_hi_hi,hi_hi_hi_hi_lo,hi_hi_hi_lo_hi,hi_hi_hi_lo_lo,hi_hi_lo_hi_hi,hi_hi_lo_hi_lo,
    hi_hi_lo_lo,hi_lo}; // @[Cat.scala 30:58]
  wire  hi_hi_hi_hi_hi_1 = reversed[62]; // @[DES_FSM.scala 173:23]
  wire  hi_hi_hi_hi_lo_1 = reversed[54]; // @[DES_FSM.scala 173:36]
  wire  hi_hi_hi_lo_hi_1 = reversed[46]; // @[DES_FSM.scala 173:49]
  wire  hi_hi_hi_lo_lo_1 = reversed[38]; // @[DES_FSM.scala 173:62]
  wire  hi_hi_lo_hi_hi_1 = reversed[30]; // @[DES_FSM.scala 173:75]
  wire  hi_hi_lo_hi_lo_1 = reversed[22]; // @[DES_FSM.scala 173:88]
  wire  hi_hi_lo_lo_1 = reversed[14]; // @[DES_FSM.scala 173:101]
  wire  hi_lo_hi_hi_hi_1 = reversed[6]; // @[DES_FSM.scala 174:13]
  wire  hi_lo_hi_hi_lo_1 = reversed[61]; // @[DES_FSM.scala 174:25]
  wire  hi_lo_hi_lo_hi_1 = reversed[53]; // @[DES_FSM.scala 174:38]
  wire  hi_lo_hi_lo_lo_1 = reversed[45]; // @[DES_FSM.scala 174:51]
  wire  hi_lo_lo_hi_hi_1 = reversed[37]; // @[DES_FSM.scala 174:64]
  wire  hi_lo_lo_hi_lo_1 = reversed[29]; // @[DES_FSM.scala 174:77]
  wire  hi_lo_lo_lo_1 = reversed[21]; // @[DES_FSM.scala 174:90]
  wire  lo_hi_hi_hi_hi_1 = reversed[13]; // @[DES_FSM.scala 175:13]
  wire  lo_hi_hi_hi_lo_1 = reversed[5]; // @[DES_FSM.scala 175:26]
  wire  lo_hi_hi_lo_hi_1 = reversed[60]; // @[DES_FSM.scala 175:38]
  wire  lo_hi_hi_lo_lo_1 = reversed[52]; // @[DES_FSM.scala 175:51]
  wire  lo_hi_lo_hi_hi_1 = reversed[44]; // @[DES_FSM.scala 175:64]
  wire  lo_hi_lo_hi_lo_1 = reversed[36]; // @[DES_FSM.scala 175:77]
  wire  lo_hi_lo_lo_1 = reversed[28]; // @[DES_FSM.scala 175:90]
  wire  lo_lo_hi_hi_hi_1 = reversed[20]; // @[DES_FSM.scala 176:13]
  wire  lo_lo_hi_hi_lo_1 = reversed[12]; // @[DES_FSM.scala 176:26]
  wire  lo_lo_hi_lo_hi_1 = reversed[4]; // @[DES_FSM.scala 176:39]
  wire  lo_lo_hi_lo_lo_1 = reversed[27]; // @[DES_FSM.scala 176:51]
  wire  lo_lo_lo_hi_hi_1 = reversed[19]; // @[DES_FSM.scala 176:64]
  wire  lo_lo_lo_hi_lo_1 = reversed[11]; // @[DES_FSM.scala 176:77]
  wire  lo_lo_lo_lo_1 = reversed[3]; // @[DES_FSM.scala 176:90]
  wire [6:0] lo_lo_1 = {lo_lo_hi_hi_hi_1,lo_lo_hi_hi_lo_1,lo_lo_hi_lo_hi_1,lo_lo_hi_lo_lo_1,lo_lo_lo_hi_hi_1,
    lo_lo_lo_hi_lo_1,lo_lo_lo_lo_1}; // @[Cat.scala 30:58]
  wire [13:0] lo_1 = {lo_hi_hi_hi_hi_1,lo_hi_hi_hi_lo_1,lo_hi_hi_lo_hi_1,lo_hi_hi_lo_lo_1,lo_hi_lo_hi_hi_1,
    lo_hi_lo_hi_lo_1,lo_hi_lo_lo_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [6:0] hi_lo_1 = {hi_lo_hi_hi_hi_1,hi_lo_hi_hi_lo_1,hi_lo_hi_lo_hi_1,hi_lo_hi_lo_lo_1,hi_lo_lo_hi_hi_1,
    hi_lo_lo_hi_lo_1,hi_lo_lo_lo_1}; // @[Cat.scala 30:58]
  wire [13:0] hi_1 = {hi_hi_hi_hi_hi_1,hi_hi_hi_hi_lo_1,hi_hi_hi_lo_hi_1,hi_hi_hi_lo_lo_1,hi_hi_lo_hi_hi_1,
    hi_hi_lo_hi_lo_1,hi_hi_lo_lo_1,hi_lo_1}; // @[Cat.scala 30:58]
  assign io_C = {hi,lo}; // @[Cat.scala 30:58]
  assign io_D = {hi_1,lo_1}; // @[Cat.scala 30:58]
endmodule
module DES_InitialPermutation(
  input  [63:0] io_text,
  input  [63:0] io_key,
  output [31:0] io_out_L,
  output [31:0] io_out_R,
  output [27:0] io_out_C,
  output [27:0] io_out_D
);
  wire [63:0] IP_io_text; // @[DES_FSM.scala 82:18]
  wire [31:0] IP_io_L; // @[DES_FSM.scala 82:18]
  wire [31:0] IP_io_R; // @[DES_FSM.scala 82:18]
  wire [63:0] PC_1_io_key; // @[DES_FSM.scala 87:20]
  wire [27:0] PC_1_io_C; // @[DES_FSM.scala 87:20]
  wire [27:0] PC_1_io_D; // @[DES_FSM.scala 87:20]
  IP IP ( // @[DES_FSM.scala 82:18]
    .io_text(IP_io_text),
    .io_L(IP_io_L),
    .io_R(IP_io_R)
  );
  PC_1 PC_1 ( // @[DES_FSM.scala 87:20]
    .io_key(PC_1_io_key),
    .io_C(PC_1_io_C),
    .io_D(PC_1_io_D)
  );
  assign io_out_L = IP_io_L; // @[DES_FSM.scala 84:12]
  assign io_out_R = IP_io_R; // @[DES_FSM.scala 85:12]
  assign io_out_C = PC_1_io_C; // @[DES_FSM.scala 89:12]
  assign io_out_D = PC_1_io_D; // @[DES_FSM.scala 90:12]
  assign IP_io_text = io_text; // @[DES_FSM.scala 83:11]
  assign PC_1_io_key = io_key; // @[DES_FSM.scala 88:12]
endmodule
module DES_FinalPermutation(
  input  [31:0] io_L,
  input  [31:0] io_R,
  output [63:0] io_out
);
  wire [63:0] _T = {io_R,io_L}; // @[Cat.scala 30:58]
  wire [63:0] _T_4 = {{32'd0}, _T[63:32]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_6 = {_T[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_8 = _T_6 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_9 = _T_4 | _T_8; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_0 = {{16'd0}, _T_9[63:16]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_14 = _GEN_0 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_16 = {_T_9[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_18 = _T_16 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_19 = _T_14 | _T_18; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_1 = {{8'd0}, _T_19[63:8]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_24 = _GEN_1 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_26 = {_T_19[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_28 = _T_26 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  wire [63:0] _T_29 = _T_24 | _T_28; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_2 = {{4'd0}, _T_29[63:4]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_34 = _GEN_2 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  wire [63:0] _T_36 = {_T_29[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_38 = _T_36 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  wire [63:0] _T_39 = _T_34 | _T_38; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_3 = {{2'd0}, _T_39[63:2]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_44 = _GEN_3 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  wire [63:0] _T_46 = {_T_39[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_48 = _T_46 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  wire [63:0] _T_49 = _T_44 | _T_48; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_4 = {{1'd0}, _T_49[63:1]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_54 = _GEN_4 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  wire [63:0] _T_56 = {_T_49[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_58 = _T_56 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  wire [63:0] concat = _T_54 | _T_58; // @[Bitwise.scala 103:39]
  wire  hi_hi_hi_hi_hi_hi = concat[39]; // @[DES_FSM.scala 127:23]
  wire  hi_hi_hi_hi_hi_lo = concat[7]; // @[DES_FSM.scala 127:34]
  wire  hi_hi_hi_hi_lo_hi = concat[47]; // @[DES_FSM.scala 127:44]
  wire  hi_hi_hi_hi_lo_lo = concat[15]; // @[DES_FSM.scala 127:55]
  wire  hi_hi_hi_lo_hi_hi = concat[55]; // @[DES_FSM.scala 127:66]
  wire  hi_hi_hi_lo_hi_lo = concat[23]; // @[DES_FSM.scala 127:77]
  wire  hi_hi_hi_lo_lo_hi = concat[63]; // @[DES_FSM.scala 127:88]
  wire  hi_hi_hi_lo_lo_lo = concat[31]; // @[DES_FSM.scala 127:99]
  wire  hi_hi_lo_hi_hi_hi = concat[38]; // @[DES_FSM.scala 128:11]
  wire  hi_hi_lo_hi_hi_lo = concat[6]; // @[DES_FSM.scala 128:22]
  wire  hi_hi_lo_hi_lo_hi = concat[46]; // @[DES_FSM.scala 128:32]
  wire  hi_hi_lo_hi_lo_lo = concat[14]; // @[DES_FSM.scala 128:43]
  wire  hi_hi_lo_lo_hi_hi = concat[54]; // @[DES_FSM.scala 128:54]
  wire  hi_hi_lo_lo_hi_lo = concat[22]; // @[DES_FSM.scala 128:65]
  wire  hi_hi_lo_lo_lo_hi = concat[62]; // @[DES_FSM.scala 128:76]
  wire  hi_hi_lo_lo_lo_lo = concat[30]; // @[DES_FSM.scala 128:87]
  wire  hi_lo_hi_hi_hi_hi = concat[37]; // @[DES_FSM.scala 129:11]
  wire  hi_lo_hi_hi_hi_lo = concat[5]; // @[DES_FSM.scala 129:22]
  wire  hi_lo_hi_hi_lo_hi = concat[45]; // @[DES_FSM.scala 129:32]
  wire  hi_lo_hi_hi_lo_lo = concat[13]; // @[DES_FSM.scala 129:43]
  wire  hi_lo_hi_lo_hi_hi = concat[53]; // @[DES_FSM.scala 129:54]
  wire  hi_lo_hi_lo_hi_lo = concat[21]; // @[DES_FSM.scala 129:65]
  wire  hi_lo_hi_lo_lo_hi = concat[61]; // @[DES_FSM.scala 129:76]
  wire  hi_lo_hi_lo_lo_lo = concat[29]; // @[DES_FSM.scala 129:87]
  wire  hi_lo_lo_hi_hi_hi = concat[36]; // @[DES_FSM.scala 130:11]
  wire  hi_lo_lo_hi_hi_lo = concat[4]; // @[DES_FSM.scala 130:22]
  wire  hi_lo_lo_hi_lo_hi = concat[44]; // @[DES_FSM.scala 130:32]
  wire  hi_lo_lo_hi_lo_lo = concat[12]; // @[DES_FSM.scala 130:43]
  wire  hi_lo_lo_lo_hi_hi = concat[52]; // @[DES_FSM.scala 130:54]
  wire  hi_lo_lo_lo_hi_lo = concat[20]; // @[DES_FSM.scala 130:65]
  wire  hi_lo_lo_lo_lo_hi = concat[60]; // @[DES_FSM.scala 130:76]
  wire  hi_lo_lo_lo_lo_lo = concat[28]; // @[DES_FSM.scala 130:87]
  wire  lo_hi_hi_hi_hi_hi = concat[35]; // @[DES_FSM.scala 131:11]
  wire  lo_hi_hi_hi_hi_lo = concat[3]; // @[DES_FSM.scala 131:22]
  wire  lo_hi_hi_hi_lo_hi = concat[43]; // @[DES_FSM.scala 131:32]
  wire  lo_hi_hi_hi_lo_lo = concat[11]; // @[DES_FSM.scala 131:43]
  wire  lo_hi_hi_lo_hi_hi = concat[51]; // @[DES_FSM.scala 131:54]
  wire  lo_hi_hi_lo_hi_lo = concat[19]; // @[DES_FSM.scala 131:65]
  wire  lo_hi_hi_lo_lo_hi = concat[59]; // @[DES_FSM.scala 131:76]
  wire  lo_hi_hi_lo_lo_lo = concat[27]; // @[DES_FSM.scala 131:87]
  wire  lo_hi_lo_hi_hi_hi = concat[34]; // @[DES_FSM.scala 132:11]
  wire  lo_hi_lo_hi_hi_lo = concat[2]; // @[DES_FSM.scala 132:22]
  wire  lo_hi_lo_hi_lo_hi = concat[42]; // @[DES_FSM.scala 132:32]
  wire  lo_hi_lo_hi_lo_lo = concat[10]; // @[DES_FSM.scala 132:43]
  wire  lo_hi_lo_lo_hi_hi = concat[50]; // @[DES_FSM.scala 132:54]
  wire  lo_hi_lo_lo_hi_lo = concat[18]; // @[DES_FSM.scala 132:65]
  wire  lo_hi_lo_lo_lo_hi = concat[58]; // @[DES_FSM.scala 132:76]
  wire  lo_hi_lo_lo_lo_lo = concat[26]; // @[DES_FSM.scala 132:87]
  wire  lo_lo_hi_hi_hi_hi = concat[33]; // @[DES_FSM.scala 133:11]
  wire  lo_lo_hi_hi_hi_lo = concat[1]; // @[DES_FSM.scala 133:22]
  wire  lo_lo_hi_hi_lo_hi = concat[41]; // @[DES_FSM.scala 133:32]
  wire  lo_lo_hi_hi_lo_lo = concat[9]; // @[DES_FSM.scala 133:43]
  wire  lo_lo_hi_lo_hi_hi = concat[49]; // @[DES_FSM.scala 133:53]
  wire  lo_lo_hi_lo_hi_lo = concat[17]; // @[DES_FSM.scala 133:64]
  wire  lo_lo_hi_lo_lo_hi = concat[57]; // @[DES_FSM.scala 133:75]
  wire  lo_lo_hi_lo_lo_lo = concat[25]; // @[DES_FSM.scala 133:86]
  wire  lo_lo_lo_hi_hi_hi = concat[32]; // @[DES_FSM.scala 134:11]
  wire  lo_lo_lo_hi_hi_lo = concat[0]; // @[DES_FSM.scala 134:22]
  wire  lo_lo_lo_hi_lo_hi = concat[40]; // @[DES_FSM.scala 134:32]
  wire  lo_lo_lo_hi_lo_lo = concat[8]; // @[DES_FSM.scala 134:43]
  wire  lo_lo_lo_lo_hi_hi = concat[48]; // @[DES_FSM.scala 134:53]
  wire  lo_lo_lo_lo_hi_lo = concat[16]; // @[DES_FSM.scala 134:64]
  wire  lo_lo_lo_lo_lo_hi = concat[56]; // @[DES_FSM.scala 134:75]
  wire  lo_lo_lo_lo_lo_lo = concat[24]; // @[DES_FSM.scala 134:86]
  wire [7:0] lo_lo_lo = {lo_lo_lo_hi_hi_hi,lo_lo_lo_hi_hi_lo,lo_lo_lo_hi_lo_hi,lo_lo_lo_hi_lo_lo,lo_lo_lo_lo_hi_hi,
    lo_lo_lo_lo_hi_lo,lo_lo_lo_lo_lo_hi,lo_lo_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [15:0] lo_lo = {lo_lo_hi_hi_hi_hi,lo_lo_hi_hi_hi_lo,lo_lo_hi_hi_lo_hi,lo_lo_hi_hi_lo_lo,lo_lo_hi_lo_hi_hi,
    lo_lo_hi_lo_hi_lo,lo_lo_hi_lo_lo_hi,lo_lo_hi_lo_lo_lo,lo_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] lo_hi_lo = {lo_hi_lo_hi_hi_hi,lo_hi_lo_hi_hi_lo,lo_hi_lo_hi_lo_hi,lo_hi_lo_hi_lo_lo,lo_hi_lo_lo_hi_hi,
    lo_hi_lo_lo_hi_lo,lo_hi_lo_lo_lo_hi,lo_hi_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [31:0] lo = {lo_hi_hi_hi_hi_hi,lo_hi_hi_hi_hi_lo,lo_hi_hi_hi_lo_hi,lo_hi_hi_hi_lo_lo,lo_hi_hi_lo_hi_hi,
    lo_hi_hi_lo_hi_lo,lo_hi_hi_lo_lo_hi,lo_hi_hi_lo_lo_lo,lo_hi_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo_lo = {hi_lo_lo_hi_hi_hi,hi_lo_lo_hi_hi_lo,hi_lo_lo_hi_lo_hi,hi_lo_lo_hi_lo_lo,hi_lo_lo_lo_hi_hi,
    hi_lo_lo_lo_hi_lo,hi_lo_lo_lo_lo_hi,hi_lo_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [15:0] hi_lo = {hi_lo_hi_hi_hi_hi,hi_lo_hi_hi_hi_lo,hi_lo_hi_hi_lo_hi,hi_lo_hi_hi_lo_lo,hi_lo_hi_lo_hi_hi,
    hi_lo_hi_lo_hi_lo,hi_lo_hi_lo_lo_hi,hi_lo_hi_lo_lo_lo,hi_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_hi_lo = {hi_hi_lo_hi_hi_hi,hi_hi_lo_hi_hi_lo,hi_hi_lo_hi_lo_hi,hi_hi_lo_hi_lo_lo,hi_hi_lo_lo_hi_hi,
    hi_hi_lo_lo_hi_lo,hi_hi_lo_lo_lo_hi,hi_hi_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [31:0] hi = {hi_hi_hi_hi_hi_hi,hi_hi_hi_hi_hi_lo,hi_hi_hi_hi_lo_hi,hi_hi_hi_hi_lo_lo,hi_hi_hi_lo_hi_hi,
    hi_hi_hi_lo_hi_lo,hi_hi_hi_lo_lo_hi,hi_hi_hi_lo_lo_lo,hi_hi_lo,hi_lo}; // @[Cat.scala 30:58]
  assign io_out = {hi,lo}; // @[Cat.scala 30:58]
endmodule
module DES_keys(
  input  [4:0]  io_round,
  input  [27:0] io_C,
  input  [27:0] io_D,
  output [27:0] io_C_next,
  output [27:0] io_D_next,
  output [47:0] io_K
);
  wire [5:0] r = {{1'd0}, io_round}; // @[DES_FSM.scala 189:15 DES_FSM.scala 193:7]
  wire  _T = 6'h0 == r; // @[Conditional.scala 37:30]
  wire  _T_1 = 6'h1 == r; // @[Conditional.scala 37:30]
  wire  _T_2 = 6'h2 == r; // @[Conditional.scala 37:30]
  wire  _T_3 = 6'h3 == r; // @[Conditional.scala 37:30]
  wire  _T_4 = 6'h4 == r; // @[Conditional.scala 37:30]
  wire  _T_5 = 6'h5 == r; // @[Conditional.scala 37:30]
  wire  _T_6 = 6'h6 == r; // @[Conditional.scala 37:30]
  wire  _T_7 = 6'h7 == r; // @[Conditional.scala 37:30]
  wire  _T_8 = 6'h8 == r; // @[Conditional.scala 37:30]
  wire  _T_9 = 6'h9 == r; // @[Conditional.scala 37:30]
  wire  _T_10 = 6'ha == r; // @[Conditional.scala 37:30]
  wire  _T_11 = 6'hb == r; // @[Conditional.scala 37:30]
  wire  _T_12 = 6'hc == r; // @[Conditional.scala 37:30]
  wire  _T_13 = 6'hd == r; // @[Conditional.scala 37:30]
  wire  _T_14 = 6'he == r; // @[Conditional.scala 37:30]
  wire  _T_15 = 6'hf == r; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_2 = _T_14 ? 2'h2 : {{1'd0}, _T_15}; // @[Conditional.scala 39:67 DES_FSM.scala 243:9]
  wire [1:0] _GEN_3 = _T_13 ? 2'h2 : _GEN_2; // @[Conditional.scala 39:67 DES_FSM.scala 240:9]
  wire [1:0] _GEN_4 = _T_12 ? 2'h2 : _GEN_3; // @[Conditional.scala 39:67 DES_FSM.scala 237:9]
  wire [1:0] _GEN_5 = _T_11 ? 2'h2 : _GEN_4; // @[Conditional.scala 39:67 DES_FSM.scala 234:9]
  wire [1:0] _GEN_6 = _T_10 ? 2'h2 : _GEN_5; // @[Conditional.scala 39:67 DES_FSM.scala 231:9]
  wire [1:0] _GEN_7 = _T_9 ? 2'h2 : _GEN_6; // @[Conditional.scala 39:67 DES_FSM.scala 228:9]
  wire [1:0] _GEN_8 = _T_8 ? 2'h1 : _GEN_7; // @[Conditional.scala 39:67 DES_FSM.scala 225:9]
  wire [1:0] _GEN_9 = _T_7 ? 2'h2 : _GEN_8; // @[Conditional.scala 39:67 DES_FSM.scala 222:9]
  wire [1:0] _GEN_10 = _T_6 ? 2'h2 : _GEN_9; // @[Conditional.scala 39:67 DES_FSM.scala 219:9]
  wire [1:0] _GEN_11 = _T_5 ? 2'h2 : _GEN_10; // @[Conditional.scala 39:67 DES_FSM.scala 216:9]
  wire [1:0] _GEN_12 = _T_4 ? 2'h2 : _GEN_11; // @[Conditional.scala 39:67 DES_FSM.scala 213:9]
  wire [1:0] _GEN_13 = _T_3 ? 2'h2 : _GEN_12; // @[Conditional.scala 39:67 DES_FSM.scala 210:9]
  wire [1:0] _GEN_14 = _T_2 ? 2'h2 : _GEN_13; // @[Conditional.scala 39:67 DES_FSM.scala 207:9]
  wire [1:0] _GEN_15 = _T_1 ? 2'h1 : _GEN_14; // @[Conditional.scala 39:67 DES_FSM.scala 204:9]
  wire [1:0] s = _T ? 2'h1 : _GEN_15; // @[Conditional.scala 40:58 DES_FSM.scala 201:9]
  wire [26:0] hi = io_C[26:0]; // @[DES_FSM.scala 259:28]
  wire  lo = io_C[27]; // @[DES_FSM.scala 259:39]
  wire [27:0] _T_18 = {hi,lo}; // @[Cat.scala 30:58]
  wire [26:0] hi_1 = io_D[26:0]; // @[DES_FSM.scala 260:28]
  wire  lo_1 = io_D[27]; // @[DES_FSM.scala 260:39]
  wire [27:0] _T_19 = {hi_1,lo_1}; // @[Cat.scala 30:58]
  wire [25:0] hi_2 = io_C[25:0]; // @[DES_FSM.scala 262:28]
  wire [1:0] lo_2 = io_C[27:26]; // @[DES_FSM.scala 262:39]
  wire [27:0] _T_20 = {hi_2,lo_2}; // @[Cat.scala 30:58]
  wire [25:0] hi_3 = io_D[25:0]; // @[DES_FSM.scala 263:28]
  wire [1:0] lo_3 = io_D[27:26]; // @[DES_FSM.scala 263:39]
  wire [27:0] _T_21 = {hi_3,lo_3}; // @[Cat.scala 30:58]
  wire [27:0] C_rotated = s == 2'h1 ? _T_18 : _T_20; // @[DES_FSM.scala 258:21 DES_FSM.scala 259:17 DES_FSM.scala 262:17]
  wire [27:0] D_rotated = s == 2'h1 ? _T_19 : _T_21; // @[DES_FSM.scala 258:21 DES_FSM.scala 260:17 DES_FSM.scala 263:17]
  wire [55:0] _T_22 = {C_rotated,D_rotated}; // @[Cat.scala 30:58]
  wire [31:0] _T_27 = {{16'd0}, _T_22[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_29 = {_T_22[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_31 = _T_29 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_32 = _T_27 | _T_31; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_19 = {{8'd0}, _T_32[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_37 = _GEN_19 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_39 = {_T_32[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_41 = _T_39 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_20 = {{4'd0}, _T_42[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_47 = _GEN_20 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_49 = {_T_42[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_51 = _T_49 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_52 = _T_47 | _T_51; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_21 = {{2'd0}, _T_52[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_57 = _GEN_21 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_59 = {_T_52[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_61 = _T_59 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_62 = _T_57 | _T_61; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_22 = {{1'd0}, _T_62[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_67 = _GEN_22 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_69 = {_T_62[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_71 = _T_69 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] hi_4 = _T_67 | _T_71; // @[Bitwise.scala 103:39]
  wire [15:0] _T_77 = {{8'd0}, _T_22[47:40]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_79 = {_T_22[39:32], 8'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_81 = _T_79 & 16'hff00; // @[Bitwise.scala 103:75]
  wire [15:0] _T_82 = _T_77 | _T_81; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_23 = {{4'd0}, _T_82[15:4]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_87 = _GEN_23 & 16'hf0f; // @[Bitwise.scala 103:31]
  wire [15:0] _T_89 = {_T_82[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_91 = _T_89 & 16'hf0f0; // @[Bitwise.scala 103:75]
  wire [15:0] _T_92 = _T_87 | _T_91; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_24 = {{2'd0}, _T_92[15:2]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_97 = _GEN_24 & 16'h3333; // @[Bitwise.scala 103:31]
  wire [15:0] _T_99 = {_T_92[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_101 = _T_99 & 16'hcccc; // @[Bitwise.scala 103:75]
  wire [15:0] _T_102 = _T_97 | _T_101; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_25 = {{1'd0}, _T_102[15:1]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_107 = _GEN_25 & 16'h5555; // @[Bitwise.scala 103:31]
  wire [15:0] _T_109 = {_T_102[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_111 = _T_109 & 16'haaaa; // @[Bitwise.scala 103:75]
  wire [15:0] hi_5 = _T_107 | _T_111; // @[Bitwise.scala 103:39]
  wire [7:0] _T_116 = {{4'd0}, _T_22[55:52]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_118 = {_T_22[51:48], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_120 = _T_118 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_121 = _T_116 | _T_120; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_26 = {{2'd0}, _T_121[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_126 = _GEN_26 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_128 = {_T_121[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_130 = _T_128 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_131 = _T_126 | _T_130; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_27 = {{1'd0}, _T_131[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_136 = _GEN_27 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_138 = {_T_131[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_140 = _T_138 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] lo_4 = _T_136 | _T_140; // @[Bitwise.scala 103:39]
  wire [55:0] concat = {hi_4,hi_5,lo_4}; // @[Cat.scala 30:58]
  wire  hi_hi_hi_hi_hi_hi = concat[13]; // @[DES_FSM.scala 283:21]
  wire  hi_hi_hi_hi_hi_lo = concat[16]; // @[DES_FSM.scala 283:32]
  wire  hi_hi_hi_hi_lo = concat[10]; // @[DES_FSM.scala 283:43]
  wire  hi_hi_hi_lo_hi_hi = concat[23]; // @[DES_FSM.scala 283:54]
  wire  hi_hi_hi_lo_hi_lo = concat[0]; // @[DES_FSM.scala 283:65]
  wire  hi_hi_hi_lo_lo = concat[4]; // @[DES_FSM.scala 283:75]
  wire  hi_hi_lo_hi_hi_hi = concat[2]; // @[DES_FSM.scala 284:11]
  wire  hi_hi_lo_hi_hi_lo = concat[27]; // @[DES_FSM.scala 284:21]
  wire  hi_hi_lo_hi_lo = concat[14]; // @[DES_FSM.scala 284:32]
  wire  hi_hi_lo_lo_hi_hi = concat[5]; // @[DES_FSM.scala 284:43]
  wire  hi_hi_lo_lo_hi_lo = concat[20]; // @[DES_FSM.scala 284:53]
  wire  hi_hi_lo_lo_lo = concat[9]; // @[DES_FSM.scala 284:64]
  wire  hi_lo_hi_hi_hi_hi = concat[22]; // @[DES_FSM.scala 285:11]
  wire  hi_lo_hi_hi_hi_lo = concat[18]; // @[DES_FSM.scala 285:22]
  wire  hi_lo_hi_hi_lo = concat[11]; // @[DES_FSM.scala 285:33]
  wire  hi_lo_hi_lo_hi_hi = concat[3]; // @[DES_FSM.scala 285:44]
  wire  hi_lo_hi_lo_hi_lo = concat[25]; // @[DES_FSM.scala 285:54]
  wire  hi_lo_hi_lo_lo = concat[7]; // @[DES_FSM.scala 285:65]
  wire  hi_lo_lo_hi_hi_hi = concat[15]; // @[DES_FSM.scala 286:11]
  wire  hi_lo_lo_hi_hi_lo = concat[6]; // @[DES_FSM.scala 286:22]
  wire  hi_lo_lo_hi_lo = concat[26]; // @[DES_FSM.scala 286:32]
  wire  hi_lo_lo_lo_hi_hi = concat[19]; // @[DES_FSM.scala 286:43]
  wire  hi_lo_lo_lo_hi_lo = concat[12]; // @[DES_FSM.scala 286:54]
  wire  hi_lo_lo_lo_lo = concat[1]; // @[DES_FSM.scala 286:65]
  wire  lo_hi_hi_hi_hi_hi = concat[40]; // @[DES_FSM.scala 287:11]
  wire  lo_hi_hi_hi_hi_lo = concat[51]; // @[DES_FSM.scala 287:22]
  wire  lo_hi_hi_hi_lo = concat[30]; // @[DES_FSM.scala 287:33]
  wire  lo_hi_hi_lo_hi_hi = concat[36]; // @[DES_FSM.scala 287:44]
  wire  lo_hi_hi_lo_hi_lo = concat[46]; // @[DES_FSM.scala 287:55]
  wire  lo_hi_hi_lo_lo = concat[54]; // @[DES_FSM.scala 287:66]
  wire  lo_hi_lo_hi_hi_hi = concat[29]; // @[DES_FSM.scala 288:11]
  wire  lo_hi_lo_hi_hi_lo = concat[39]; // @[DES_FSM.scala 288:22]
  wire  lo_hi_lo_hi_lo = concat[50]; // @[DES_FSM.scala 288:33]
  wire  lo_hi_lo_lo_hi_hi = concat[44]; // @[DES_FSM.scala 288:44]
  wire  lo_hi_lo_lo_hi_lo = concat[32]; // @[DES_FSM.scala 288:55]
  wire  lo_hi_lo_lo_lo = concat[47]; // @[DES_FSM.scala 288:66]
  wire  lo_lo_hi_hi_hi_hi = concat[43]; // @[DES_FSM.scala 289:11]
  wire  lo_lo_hi_hi_hi_lo = concat[48]; // @[DES_FSM.scala 289:22]
  wire  lo_lo_hi_hi_lo = concat[38]; // @[DES_FSM.scala 289:33]
  wire  lo_lo_hi_lo_hi_hi = concat[55]; // @[DES_FSM.scala 289:44]
  wire  lo_lo_hi_lo_hi_lo = concat[33]; // @[DES_FSM.scala 289:55]
  wire  lo_lo_hi_lo_lo = concat[52]; // @[DES_FSM.scala 289:66]
  wire  lo_lo_lo_hi_hi_hi = concat[45]; // @[DES_FSM.scala 290:11]
  wire  lo_lo_lo_hi_hi_lo = concat[41]; // @[DES_FSM.scala 290:22]
  wire  lo_lo_lo_hi_lo = concat[49]; // @[DES_FSM.scala 290:33]
  wire  lo_lo_lo_lo_hi_hi = concat[35]; // @[DES_FSM.scala 290:44]
  wire  lo_lo_lo_lo_hi_lo = concat[28]; // @[DES_FSM.scala 290:55]
  wire  lo_lo_lo_lo_lo = concat[31]; // @[DES_FSM.scala 290:66]
  wire [5:0] lo_lo_lo = {lo_lo_lo_hi_hi_hi,lo_lo_lo_hi_hi_lo,lo_lo_lo_hi_lo,lo_lo_lo_lo_hi_hi,lo_lo_lo_lo_hi_lo,
    lo_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [11:0] lo_lo = {lo_lo_hi_hi_hi_hi,lo_lo_hi_hi_hi_lo,lo_lo_hi_hi_lo,lo_lo_hi_lo_hi_hi,lo_lo_hi_lo_hi_lo,
    lo_lo_hi_lo_lo,lo_lo_lo}; // @[Cat.scala 30:58]
  wire [5:0] lo_hi_lo = {lo_hi_lo_hi_hi_hi,lo_hi_lo_hi_hi_lo,lo_hi_lo_hi_lo,lo_hi_lo_lo_hi_hi,lo_hi_lo_lo_hi_lo,
    lo_hi_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [23:0] lo_6 = {lo_hi_hi_hi_hi_hi,lo_hi_hi_hi_hi_lo,lo_hi_hi_hi_lo,lo_hi_hi_lo_hi_hi,lo_hi_hi_lo_hi_lo,
    lo_hi_hi_lo_lo,lo_hi_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [5:0] hi_lo_lo = {hi_lo_lo_hi_hi_hi,hi_lo_lo_hi_hi_lo,hi_lo_lo_hi_lo,hi_lo_lo_lo_hi_hi,hi_lo_lo_lo_hi_lo,
    hi_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [11:0] hi_lo = {hi_lo_hi_hi_hi_hi,hi_lo_hi_hi_hi_lo,hi_lo_hi_hi_lo,hi_lo_hi_lo_hi_hi,hi_lo_hi_lo_hi_lo,
    hi_lo_hi_lo_lo,hi_lo_lo}; // @[Cat.scala 30:58]
  wire [5:0] hi_hi_lo = {hi_hi_lo_hi_hi_hi,hi_hi_lo_hi_hi_lo,hi_hi_lo_hi_lo,hi_hi_lo_lo_hi_hi,hi_hi_lo_lo_hi_lo,
    hi_hi_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [23:0] hi_6 = {hi_hi_hi_hi_hi_hi,hi_hi_hi_hi_hi_lo,hi_hi_hi_hi_lo,hi_hi_hi_lo_hi_hi,hi_hi_hi_lo_hi_lo,
    hi_hi_hi_lo_lo,hi_hi_lo,hi_lo}; // @[Cat.scala 30:58]
  assign io_C_next = s == 2'h1 ? _T_18 : _T_20; // @[DES_FSM.scala 258:21 DES_FSM.scala 259:17 DES_FSM.scala 262:17]
  assign io_D_next = s == 2'h1 ? _T_19 : _T_21; // @[DES_FSM.scala 258:21 DES_FSM.scala 260:17 DES_FSM.scala 263:17]
  assign io_K = {hi_6,lo_6}; // @[Cat.scala 30:58]
endmodule
module DES_E(
  input  [31:0] io_R,
  output [47:0] io_E
);
  wire [31:0] _T_3 = {{16'd0}, io_R[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_5 = {io_R[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_7 = _T_5 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_8 = _T_3 | _T_7; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_0 = {{8'd0}, _T_8[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_13 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_15 = {_T_8[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_17 = _T_15 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_18 = _T_13 | _T_17; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1 = {{4'd0}, _T_18[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_23 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_25 = {_T_18[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_27 = _T_25 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_28 = _T_23 | _T_27; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_2 = {{2'd0}, _T_28[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_33 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_35 = {_T_28[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_37 = _T_35 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_38 = _T_33 | _T_37; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3 = {{1'd0}, _T_38[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_43 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_45 = {_T_38[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_47 = _T_45 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] reversed = _T_43 | _T_47; // @[Bitwise.scala 103:39]
  wire  hi_hi_hi_hi_hi_hi = reversed[31]; // @[DES_FSM.scala 494:23]
  wire  hi_hi_hi_hi_hi_lo = reversed[0]; // @[DES_FSM.scala 494:36]
  wire  hi_hi_hi_hi_lo = reversed[1]; // @[DES_FSM.scala 494:48]
  wire  hi_hi_hi_lo_hi_hi = reversed[2]; // @[DES_FSM.scala 494:60]
  wire  hi_hi_hi_lo_hi_lo = reversed[3]; // @[DES_FSM.scala 494:72]
  wire  hi_hi_hi_lo_lo = reversed[4]; // @[DES_FSM.scala 494:84]
  wire  hi_hi_lo_hi_lo = reversed[5]; // @[DES_FSM.scala 495:37]
  wire  hi_hi_lo_lo_hi_hi = reversed[6]; // @[DES_FSM.scala 495:49]
  wire  hi_hi_lo_lo_hi_lo = reversed[7]; // @[DES_FSM.scala 495:61]
  wire  hi_hi_lo_lo_lo = reversed[8]; // @[DES_FSM.scala 495:73]
  wire  hi_lo_hi_hi_lo = reversed[9]; // @[DES_FSM.scala 496:37]
  wire  hi_lo_hi_lo_hi_hi = reversed[10]; // @[DES_FSM.scala 496:49]
  wire  hi_lo_hi_lo_hi_lo = reversed[11]; // @[DES_FSM.scala 496:62]
  wire  hi_lo_hi_lo_lo = reversed[12]; // @[DES_FSM.scala 496:75]
  wire  hi_lo_lo_hi_lo = reversed[13]; // @[DES_FSM.scala 497:39]
  wire  hi_lo_lo_lo_hi_hi = reversed[14]; // @[DES_FSM.scala 497:52]
  wire  hi_lo_lo_lo_hi_lo = reversed[15]; // @[DES_FSM.scala 497:65]
  wire  hi_lo_lo_lo_lo = reversed[16]; // @[DES_FSM.scala 497:78]
  wire  lo_hi_hi_hi_lo = reversed[17]; // @[DES_FSM.scala 498:39]
  wire  lo_hi_hi_lo_hi_hi = reversed[18]; // @[DES_FSM.scala 498:52]
  wire  lo_hi_hi_lo_hi_lo = reversed[19]; // @[DES_FSM.scala 498:65]
  wire  lo_hi_hi_lo_lo = reversed[20]; // @[DES_FSM.scala 498:78]
  wire  lo_hi_lo_hi_lo = reversed[21]; // @[DES_FSM.scala 499:39]
  wire  lo_hi_lo_lo_hi_hi = reversed[22]; // @[DES_FSM.scala 499:52]
  wire  lo_hi_lo_lo_hi_lo = reversed[23]; // @[DES_FSM.scala 499:65]
  wire  lo_hi_lo_lo_lo = reversed[24]; // @[DES_FSM.scala 499:78]
  wire  lo_lo_hi_hi_lo = reversed[25]; // @[DES_FSM.scala 500:39]
  wire  lo_lo_hi_lo_hi_hi = reversed[26]; // @[DES_FSM.scala 500:52]
  wire  lo_lo_hi_lo_hi_lo = reversed[27]; // @[DES_FSM.scala 500:65]
  wire  lo_lo_hi_lo_lo = reversed[28]; // @[DES_FSM.scala 500:78]
  wire  lo_lo_lo_hi_lo = reversed[29]; // @[DES_FSM.scala 501:39]
  wire  lo_lo_lo_lo_hi_hi = reversed[30]; // @[DES_FSM.scala 501:52]
  wire [5:0] lo_lo_lo = {lo_lo_hi_lo_hi_lo,lo_lo_hi_lo_lo,lo_lo_lo_hi_lo,lo_lo_lo_lo_hi_hi,hi_hi_hi_hi_hi_hi,
    hi_hi_hi_hi_hi_lo}; // @[Cat.scala 30:58]
  wire [11:0] lo_lo = {lo_hi_lo_lo_hi_lo,lo_hi_lo_lo_lo,lo_lo_hi_hi_lo,lo_lo_hi_lo_hi_hi,lo_lo_hi_lo_hi_lo,
    lo_lo_hi_lo_lo,lo_lo_lo}; // @[Cat.scala 30:58]
  wire [5:0] lo_hi_lo = {lo_hi_hi_lo_hi_lo,lo_hi_hi_lo_lo,lo_hi_lo_hi_lo,lo_hi_lo_lo_hi_hi,lo_hi_lo_lo_hi_lo,
    lo_hi_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [23:0] lo = {hi_lo_lo_lo_hi_lo,hi_lo_lo_lo_lo,lo_hi_hi_hi_lo,lo_hi_hi_lo_hi_hi,lo_hi_hi_lo_hi_lo,lo_hi_hi_lo_lo,
    lo_hi_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [5:0] hi_lo_lo = {hi_lo_hi_lo_hi_lo,hi_lo_hi_lo_lo,hi_lo_lo_hi_lo,hi_lo_lo_lo_hi_hi,hi_lo_lo_lo_hi_lo,
    hi_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [11:0] hi_lo = {hi_hi_lo_lo_hi_lo,hi_hi_lo_lo_lo,hi_lo_hi_hi_lo,hi_lo_hi_lo_hi_hi,hi_lo_hi_lo_hi_lo,
    hi_lo_hi_lo_lo,hi_lo_lo}; // @[Cat.scala 30:58]
  wire [5:0] hi_hi_lo = {hi_hi_hi_lo_hi_lo,hi_hi_hi_lo_lo,hi_hi_lo_hi_lo,hi_hi_lo_lo_hi_hi,hi_hi_lo_lo_hi_lo,
    hi_hi_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [23:0] hi = {hi_hi_hi_hi_hi_hi,hi_hi_hi_hi_hi_lo,hi_hi_hi_hi_lo,hi_hi_hi_lo_hi_hi,hi_hi_hi_lo_hi_lo,
    hi_hi_hi_lo_lo,hi_hi_lo,hi_lo}; // @[Cat.scala 30:58]
  assign io_E = {hi,lo}; // @[Cat.scala 30:58]
endmodule
module DES_S(
  input  [47:0] io_in,
  output [31:0] io_out
);
  wire [5:0] B_7 = io_in[5:0]; // @[DES_FSM.scala 321:20]
  wire  hi = B_7[5]; // @[DES_FSM.scala 322:27]
  wire  lo = B_7[0]; // @[DES_FSM.scala 322:37]
  wire [1:0] row_7 = {hi,lo}; // @[Cat.scala 30:58]
  wire [3:0] col_7 = B_7[4:1]; // @[DES_FSM.scala 323:23]
  wire [5:0] B_6 = io_in[11:6]; // @[DES_FSM.scala 321:20]
  wire  hi_1 = B_6[5]; // @[DES_FSM.scala 322:27]
  wire  lo_1 = B_6[0]; // @[DES_FSM.scala 322:37]
  wire [1:0] row_6 = {hi_1,lo_1}; // @[Cat.scala 30:58]
  wire [3:0] col_6 = B_6[4:1]; // @[DES_FSM.scala 323:23]
  wire [5:0] B_5 = io_in[17:12]; // @[DES_FSM.scala 321:20]
  wire  hi_2 = B_5[5]; // @[DES_FSM.scala 322:27]
  wire  lo_2 = B_5[0]; // @[DES_FSM.scala 322:37]
  wire [1:0] row_5 = {hi_2,lo_2}; // @[Cat.scala 30:58]
  wire [3:0] col_5 = B_5[4:1]; // @[DES_FSM.scala 323:23]
  wire [5:0] B_4 = io_in[23:18]; // @[DES_FSM.scala 321:20]
  wire  hi_3 = B_4[5]; // @[DES_FSM.scala 322:27]
  wire  lo_3 = B_4[0]; // @[DES_FSM.scala 322:37]
  wire [1:0] row_4 = {hi_3,lo_3}; // @[Cat.scala 30:58]
  wire [3:0] col_4 = B_4[4:1]; // @[DES_FSM.scala 323:23]
  wire [5:0] B_3 = io_in[29:24]; // @[DES_FSM.scala 321:20]
  wire  hi_4 = B_3[5]; // @[DES_FSM.scala 322:27]
  wire  lo_4 = B_3[0]; // @[DES_FSM.scala 322:37]
  wire [1:0] row_3 = {hi_4,lo_4}; // @[Cat.scala 30:58]
  wire [3:0] col_3 = B_3[4:1]; // @[DES_FSM.scala 323:23]
  wire [5:0] B_2 = io_in[35:30]; // @[DES_FSM.scala 321:20]
  wire  hi_5 = B_2[5]; // @[DES_FSM.scala 322:27]
  wire  lo_5 = B_2[0]; // @[DES_FSM.scala 322:37]
  wire [1:0] row_2 = {hi_5,lo_5}; // @[Cat.scala 30:58]
  wire [3:0] col_2 = B_2[4:1]; // @[DES_FSM.scala 323:23]
  wire [5:0] B_1 = io_in[41:36]; // @[DES_FSM.scala 321:20]
  wire  hi_6 = B_1[5]; // @[DES_FSM.scala 322:27]
  wire  lo_6 = B_1[0]; // @[DES_FSM.scala 322:37]
  wire [1:0] row_1 = {hi_6,lo_6}; // @[Cat.scala 30:58]
  wire [3:0] col_1 = B_1[4:1]; // @[DES_FSM.scala 323:23]
  wire [5:0] B_0 = io_in[47:42]; // @[DES_FSM.scala 321:20]
  wire  hi_7 = B_0[5]; // @[DES_FSM.scala 322:27]
  wire  lo_7 = B_0[0]; // @[DES_FSM.scala 322:37]
  wire [1:0] row_0 = {hi_7,lo_7}; // @[Cat.scala 30:58]
  wire [3:0] col_0 = B_0[4:1]; // @[DES_FSM.scala 323:23]
  wire [3:0] _GEN_1 = 4'h0 == col_6 & 2'h1 == row_6 ? 4'hd : 4'h4; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_2 = 4'h0 == col_6 & 2'h2 == row_6 ? 4'h1 : _GEN_1; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_3 = 4'h0 == col_6 & 2'h3 == row_6 ? 4'h6 : _GEN_2; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_4 = 4'h1 == col_6 & 2'h0 == row_6 ? 4'hb : _GEN_3; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_5 = 4'h1 == col_6 & 2'h1 == row_6 ? 4'h0 : _GEN_4; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_6 = 4'h1 == col_6 & 2'h2 == row_6 ? 4'h4 : _GEN_5; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_7 = 4'h1 == col_6 & 2'h3 == row_6 ? 4'hb : _GEN_6; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_8 = 4'h2 == col_6 & 2'h0 == row_6 ? 4'h2 : _GEN_7; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_9 = 4'h2 == col_6 & 2'h1 == row_6 ? 4'hb : _GEN_8; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_10 = 4'h2 == col_6 & 2'h2 == row_6 ? 4'hb : _GEN_9; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_11 = 4'h2 == col_6 & 2'h3 == row_6 ? 4'hd : _GEN_10; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_12 = 4'h3 == col_6 & 2'h0 == row_6 ? 4'he : _GEN_11; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_13 = 4'h3 == col_6 & 2'h1 == row_6 ? 4'h7 : _GEN_12; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_14 = 4'h3 == col_6 & 2'h2 == row_6 ? 4'hd : _GEN_13; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_15 = 4'h3 == col_6 & 2'h3 == row_6 ? 4'h8 : _GEN_14; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_16 = 4'h4 == col_6 & 2'h0 == row_6 ? 4'hf : _GEN_15; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_17 = 4'h4 == col_6 & 2'h1 == row_6 ? 4'h4 : _GEN_16; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_18 = 4'h4 == col_6 & 2'h2 == row_6 ? 4'hc : _GEN_17; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_19 = 4'h4 == col_6 & 2'h3 == row_6 ? 4'h1 : _GEN_18; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_20 = 4'h5 == col_6 & 2'h0 == row_6 ? 4'h0 : _GEN_19; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_21 = 4'h5 == col_6 & 2'h1 == row_6 ? 4'h9 : _GEN_20; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_22 = 4'h5 == col_6 & 2'h2 == row_6 ? 4'h3 : _GEN_21; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_23 = 4'h5 == col_6 & 2'h3 == row_6 ? 4'h4 : _GEN_22; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_24 = 4'h6 == col_6 & 2'h0 == row_6 ? 4'h8 : _GEN_23; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_25 = 4'h6 == col_6 & 2'h1 == row_6 ? 4'h1 : _GEN_24; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_26 = 4'h6 == col_6 & 2'h2 == row_6 ? 4'h7 : _GEN_25; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_27 = 4'h6 == col_6 & 2'h3 == row_6 ? 4'ha : _GEN_26; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_28 = 4'h7 == col_6 & 2'h0 == row_6 ? 4'hd : _GEN_27; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_29 = 4'h7 == col_6 & 2'h1 == row_6 ? 4'ha : _GEN_28; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_30 = 4'h7 == col_6 & 2'h2 == row_6 ? 4'he : _GEN_29; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_31 = 4'h7 == col_6 & 2'h3 == row_6 ? 4'h7 : _GEN_30; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_32 = 4'h8 == col_6 & 2'h0 == row_6 ? 4'h3 : _GEN_31; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_33 = 4'h8 == col_6 & 2'h1 == row_6 ? 4'he : _GEN_32; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_34 = 4'h8 == col_6 & 2'h2 == row_6 ? 4'ha : _GEN_33; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_35 = 4'h8 == col_6 & 2'h3 == row_6 ? 4'h9 : _GEN_34; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_36 = 4'h9 == col_6 & 2'h0 == row_6 ? 4'hc : _GEN_35; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_37 = 4'h9 == col_6 & 2'h1 == row_6 ? 4'h3 : _GEN_36; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_38 = 4'h9 == col_6 & 2'h2 == row_6 ? 4'hf : _GEN_37; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_39 = 4'h9 == col_6 & 2'h3 == row_6 ? 4'h5 : _GEN_38; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_40 = 4'ha == col_6 & 2'h0 == row_6 ? 4'h9 : _GEN_39; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_41 = 4'ha == col_6 & 2'h1 == row_6 ? 4'h5 : _GEN_40; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_42 = 4'ha == col_6 & 2'h2 == row_6 ? 4'h6 : _GEN_41; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_43 = 4'ha == col_6 & 2'h3 == row_6 ? 4'h0 : _GEN_42; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_44 = 4'hb == col_6 & 2'h0 == row_6 ? 4'h7 : _GEN_43; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_45 = 4'hb == col_6 & 2'h1 == row_6 ? 4'hc : _GEN_44; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_46 = 4'hb == col_6 & 2'h2 == row_6 ? 4'h8 : _GEN_45; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_47 = 4'hb == col_6 & 2'h3 == row_6 ? 4'hf : _GEN_46; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_48 = 4'hc == col_6 & 2'h0 == row_6 ? 4'h5 : _GEN_47; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_49 = 4'hc == col_6 & 2'h1 == row_6 ? 4'h2 : _GEN_48; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_50 = 4'hc == col_6 & 2'h2 == row_6 ? 4'h0 : _GEN_49; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_51 = 4'hc == col_6 & 2'h3 == row_6 ? 4'he : _GEN_50; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_52 = 4'hd == col_6 & 2'h0 == row_6 ? 4'ha : _GEN_51; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_53 = 4'hd == col_6 & 2'h1 == row_6 ? 4'hf : _GEN_52; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_54 = 4'hd == col_6 & 2'h2 == row_6 ? 4'h5 : _GEN_53; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_55 = 4'hd == col_6 & 2'h3 == row_6 ? 4'h2 : _GEN_54; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_56 = 4'he == col_6 & 2'h0 == row_6 ? 4'h6 : _GEN_55; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_57 = 4'he == col_6 & 2'h1 == row_6 ? 4'h8 : _GEN_56; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_58 = 4'he == col_6 & 2'h2 == row_6 ? 4'h9 : _GEN_57; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_59 = 4'he == col_6 & 2'h3 == row_6 ? 4'h3 : _GEN_58; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_60 = 4'hf == col_6 & 2'h0 == row_6 ? 4'h1 : _GEN_59; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_61 = 4'hf == col_6 & 2'h1 == row_6 ? 4'h6 : _GEN_60; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_62 = 4'hf == col_6 & 2'h2 == row_6 ? 4'h2 : _GEN_61; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_63 = 4'hf == col_6 & 2'h3 == row_6 ? 4'hc : _GEN_62; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_65 = 4'h0 == col_7 & 2'h1 == row_7 ? 4'h1 : 4'hd; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_66 = 4'h0 == col_7 & 2'h2 == row_7 ? 4'h7 : _GEN_65; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_67 = 4'h0 == col_7 & 2'h3 == row_7 ? 4'h2 : _GEN_66; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_68 = 4'h1 == col_7 & 2'h0 == row_7 ? 4'h2 : _GEN_67; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_69 = 4'h1 == col_7 & 2'h1 == row_7 ? 4'hf : _GEN_68; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_70 = 4'h1 == col_7 & 2'h2 == row_7 ? 4'hb : _GEN_69; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_71 = 4'h1 == col_7 & 2'h3 == row_7 ? 4'h1 : _GEN_70; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_72 = 4'h2 == col_7 & 2'h0 == row_7 ? 4'h8 : _GEN_71; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_73 = 4'h2 == col_7 & 2'h1 == row_7 ? 4'hd : _GEN_72; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_74 = 4'h2 == col_7 & 2'h2 == row_7 ? 4'h4 : _GEN_73; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_75 = 4'h2 == col_7 & 2'h3 == row_7 ? 4'he : _GEN_74; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_76 = 4'h3 == col_7 & 2'h0 == row_7 ? 4'h4 : _GEN_75; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_77 = 4'h3 == col_7 & 2'h1 == row_7 ? 4'h8 : _GEN_76; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_78 = 4'h3 == col_7 & 2'h2 == row_7 ? 4'h1 : _GEN_77; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_79 = 4'h3 == col_7 & 2'h3 == row_7 ? 4'h7 : _GEN_78; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_80 = 4'h4 == col_7 & 2'h0 == row_7 ? 4'h6 : _GEN_79; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_81 = 4'h4 == col_7 & 2'h1 == row_7 ? 4'ha : _GEN_80; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_82 = 4'h4 == col_7 & 2'h2 == row_7 ? 4'h9 : _GEN_81; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_83 = 4'h4 == col_7 & 2'h3 == row_7 ? 4'h4 : _GEN_82; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_84 = 4'h5 == col_7 & 2'h0 == row_7 ? 4'hf : _GEN_83; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_85 = 4'h5 == col_7 & 2'h1 == row_7 ? 4'h3 : _GEN_84; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_86 = 4'h5 == col_7 & 2'h2 == row_7 ? 4'hc : _GEN_85; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_87 = 4'h5 == col_7 & 2'h3 == row_7 ? 4'ha : _GEN_86; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_88 = 4'h6 == col_7 & 2'h0 == row_7 ? 4'hb : _GEN_87; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_89 = 4'h6 == col_7 & 2'h1 == row_7 ? 4'h7 : _GEN_88; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_90 = 4'h6 == col_7 & 2'h2 == row_7 ? 4'he : _GEN_89; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_91 = 4'h6 == col_7 & 2'h3 == row_7 ? 4'h8 : _GEN_90; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_92 = 4'h7 == col_7 & 2'h0 == row_7 ? 4'h1 : _GEN_91; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_93 = 4'h7 == col_7 & 2'h1 == row_7 ? 4'h4 : _GEN_92; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_94 = 4'h7 == col_7 & 2'h2 == row_7 ? 4'h2 : _GEN_93; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_95 = 4'h7 == col_7 & 2'h3 == row_7 ? 4'hd : _GEN_94; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_96 = 4'h8 == col_7 & 2'h0 == row_7 ? 4'ha : _GEN_95; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_97 = 4'h8 == col_7 & 2'h1 == row_7 ? 4'hc : _GEN_96; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_98 = 4'h8 == col_7 & 2'h2 == row_7 ? 4'h0 : _GEN_97; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_99 = 4'h8 == col_7 & 2'h3 == row_7 ? 4'hf : _GEN_98; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_100 = 4'h9 == col_7 & 2'h0 == row_7 ? 4'h9 : _GEN_99; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_101 = 4'h9 == col_7 & 2'h1 == row_7 ? 4'h5 : _GEN_100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_102 = 4'h9 == col_7 & 2'h2 == row_7 ? 4'h6 : _GEN_101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_103 = 4'h9 == col_7 & 2'h3 == row_7 ? 4'hc : _GEN_102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_104 = 4'ha == col_7 & 2'h0 == row_7 ? 4'h3 : _GEN_103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_105 = 4'ha == col_7 & 2'h1 == row_7 ? 4'h6 : _GEN_104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_106 = 4'ha == col_7 & 2'h2 == row_7 ? 4'ha : _GEN_105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_107 = 4'ha == col_7 & 2'h3 == row_7 ? 4'h9 : _GEN_106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_108 = 4'hb == col_7 & 2'h0 == row_7 ? 4'he : _GEN_107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_109 = 4'hb == col_7 & 2'h1 == row_7 ? 4'hb : _GEN_108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_110 = 4'hb == col_7 & 2'h2 == row_7 ? 4'hd : _GEN_109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_111 = 4'hb == col_7 & 2'h3 == row_7 ? 4'h0 : _GEN_110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_112 = 4'hc == col_7 & 2'h0 == row_7 ? 4'h5 : _GEN_111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_113 = 4'hc == col_7 & 2'h1 == row_7 ? 4'h0 : _GEN_112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_114 = 4'hc == col_7 & 2'h2 == row_7 ? 4'hf : _GEN_113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_115 = 4'hc == col_7 & 2'h3 == row_7 ? 4'h3 : _GEN_114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_116 = 4'hd == col_7 & 2'h0 == row_7 ? 4'h0 : _GEN_115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_117 = 4'hd == col_7 & 2'h1 == row_7 ? 4'he : _GEN_116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_118 = 4'hd == col_7 & 2'h2 == row_7 ? 4'h3 : _GEN_117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_119 = 4'hd == col_7 & 2'h3 == row_7 ? 4'h5 : _GEN_118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_120 = 4'he == col_7 & 2'h0 == row_7 ? 4'hc : _GEN_119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_121 = 4'he == col_7 & 2'h1 == row_7 ? 4'h9 : _GEN_120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_122 = 4'he == col_7 & 2'h2 == row_7 ? 4'h5 : _GEN_121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_123 = 4'he == col_7 & 2'h3 == row_7 ? 4'h6 : _GEN_122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_124 = 4'hf == col_7 & 2'h0 == row_7 ? 4'h7 : _GEN_123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_125 = 4'hf == col_7 & 2'h1 == row_7 ? 4'h2 : _GEN_124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_126 = 4'hf == col_7 & 2'h2 == row_7 ? 4'h8 : _GEN_125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_127 = 4'hf == col_7 & 2'h3 == row_7 ? 4'hb : _GEN_126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_129 = 4'h0 == col_4 & 2'h1 == row_4 ? 4'he : 4'h2; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_130 = 4'h0 == col_4 & 2'h2 == row_4 ? 4'h4 : _GEN_129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_131 = 4'h0 == col_4 & 2'h3 == row_4 ? 4'hb : _GEN_130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_132 = 4'h1 == col_4 & 2'h0 == row_4 ? 4'hc : _GEN_131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_133 = 4'h1 == col_4 & 2'h1 == row_4 ? 4'hb : _GEN_132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_134 = 4'h1 == col_4 & 2'h2 == row_4 ? 4'h2 : _GEN_133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_135 = 4'h1 == col_4 & 2'h3 == row_4 ? 4'h8 : _GEN_134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_136 = 4'h2 == col_4 & 2'h0 == row_4 ? 4'h4 : _GEN_135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_137 = 4'h2 == col_4 & 2'h1 == row_4 ? 4'h2 : _GEN_136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_138 = 4'h2 == col_4 & 2'h2 == row_4 ? 4'h1 : _GEN_137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_139 = 4'h2 == col_4 & 2'h3 == row_4 ? 4'hc : _GEN_138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_140 = 4'h3 == col_4 & 2'h0 == row_4 ? 4'h1 : _GEN_139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_141 = 4'h3 == col_4 & 2'h1 == row_4 ? 4'hc : _GEN_140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_142 = 4'h3 == col_4 & 2'h2 == row_4 ? 4'hb : _GEN_141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_143 = 4'h3 == col_4 & 2'h3 == row_4 ? 4'h7 : _GEN_142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_144 = 4'h4 == col_4 & 2'h0 == row_4 ? 4'h7 : _GEN_143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_145 = 4'h4 == col_4 & 2'h1 == row_4 ? 4'h4 : _GEN_144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_146 = 4'h4 == col_4 & 2'h2 == row_4 ? 4'ha : _GEN_145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_147 = 4'h4 == col_4 & 2'h3 == row_4 ? 4'h1 : _GEN_146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_148 = 4'h5 == col_4 & 2'h0 == row_4 ? 4'ha : _GEN_147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_149 = 4'h5 == col_4 & 2'h1 == row_4 ? 4'h7 : _GEN_148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_150 = 4'h5 == col_4 & 2'h2 == row_4 ? 4'hd : _GEN_149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_151 = 4'h5 == col_4 & 2'h3 == row_4 ? 4'he : _GEN_150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_152 = 4'h6 == col_4 & 2'h0 == row_4 ? 4'hb : _GEN_151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_153 = 4'h6 == col_4 & 2'h1 == row_4 ? 4'hd : _GEN_152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_154 = 4'h6 == col_4 & 2'h2 == row_4 ? 4'h7 : _GEN_153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_155 = 4'h6 == col_4 & 2'h3 == row_4 ? 4'h2 : _GEN_154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_156 = 4'h7 == col_4 & 2'h0 == row_4 ? 4'h6 : _GEN_155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_157 = 4'h7 == col_4 & 2'h1 == row_4 ? 4'h1 : _GEN_156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_158 = 4'h7 == col_4 & 2'h2 == row_4 ? 4'h8 : _GEN_157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_159 = 4'h7 == col_4 & 2'h3 == row_4 ? 4'hd : _GEN_158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_160 = 4'h8 == col_4 & 2'h0 == row_4 ? 4'h8 : _GEN_159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_161 = 4'h8 == col_4 & 2'h1 == row_4 ? 4'h5 : _GEN_160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_162 = 4'h8 == col_4 & 2'h2 == row_4 ? 4'hf : _GEN_161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_163 = 4'h8 == col_4 & 2'h3 == row_4 ? 4'h6 : _GEN_162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_164 = 4'h9 == col_4 & 2'h0 == row_4 ? 4'h5 : _GEN_163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_165 = 4'h9 == col_4 & 2'h1 == row_4 ? 4'h0 : _GEN_164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_166 = 4'h9 == col_4 & 2'h2 == row_4 ? 4'h9 : _GEN_165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_167 = 4'h9 == col_4 & 2'h3 == row_4 ? 4'hf : _GEN_166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_168 = 4'ha == col_4 & 2'h0 == row_4 ? 4'h3 : _GEN_167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_169 = 4'ha == col_4 & 2'h1 == row_4 ? 4'hf : _GEN_168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_170 = 4'ha == col_4 & 2'h2 == row_4 ? 4'hc : _GEN_169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_171 = 4'ha == col_4 & 2'h3 == row_4 ? 4'h0 : _GEN_170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_172 = 4'hb == col_4 & 2'h0 == row_4 ? 4'hf : _GEN_171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_173 = 4'hb == col_4 & 2'h1 == row_4 ? 4'ha : _GEN_172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_174 = 4'hb == col_4 & 2'h2 == row_4 ? 4'h5 : _GEN_173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_175 = 4'hb == col_4 & 2'h3 == row_4 ? 4'h9 : _GEN_174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_176 = 4'hc == col_4 & 2'h0 == row_4 ? 4'hd : _GEN_175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_177 = 4'hc == col_4 & 2'h1 == row_4 ? 4'h3 : _GEN_176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_178 = 4'hc == col_4 & 2'h2 == row_4 ? 4'h6 : _GEN_177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_179 = 4'hc == col_4 & 2'h3 == row_4 ? 4'ha : _GEN_178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_180 = 4'hd == col_4 & 2'h0 == row_4 ? 4'h0 : _GEN_179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_181 = 4'hd == col_4 & 2'h1 == row_4 ? 4'h9 : _GEN_180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_182 = 4'hd == col_4 & 2'h2 == row_4 ? 4'h3 : _GEN_181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_183 = 4'hd == col_4 & 2'h3 == row_4 ? 4'h4 : _GEN_182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_184 = 4'he == col_4 & 2'h0 == row_4 ? 4'he : _GEN_183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_185 = 4'he == col_4 & 2'h1 == row_4 ? 4'h8 : _GEN_184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_186 = 4'he == col_4 & 2'h2 == row_4 ? 4'h0 : _GEN_185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_187 = 4'he == col_4 & 2'h3 == row_4 ? 4'h5 : _GEN_186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_188 = 4'hf == col_4 & 2'h0 == row_4 ? 4'h9 : _GEN_187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_189 = 4'hf == col_4 & 2'h1 == row_4 ? 4'h6 : _GEN_188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_190 = 4'hf == col_4 & 2'h2 == row_4 ? 4'he : _GEN_189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_191 = 4'hf == col_4 & 2'h3 == row_4 ? 4'h3 : _GEN_190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_193 = 4'h0 == col_5 & 2'h1 == row_5 ? 4'ha : 4'hc; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_194 = 4'h0 == col_5 & 2'h2 == row_5 ? 4'h9 : _GEN_193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_195 = 4'h0 == col_5 & 2'h3 == row_5 ? 4'h4 : _GEN_194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_196 = 4'h1 == col_5 & 2'h0 == row_5 ? 4'h1 : _GEN_195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_197 = 4'h1 == col_5 & 2'h1 == row_5 ? 4'hf : _GEN_196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_198 = 4'h1 == col_5 & 2'h2 == row_5 ? 4'he : _GEN_197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_199 = 4'h1 == col_5 & 2'h3 == row_5 ? 4'h3 : _GEN_198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_200 = 4'h2 == col_5 & 2'h0 == row_5 ? 4'ha : _GEN_199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_201 = 4'h2 == col_5 & 2'h1 == row_5 ? 4'h4 : _GEN_200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_202 = 4'h2 == col_5 & 2'h2 == row_5 ? 4'hf : _GEN_201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_203 = 4'h2 == col_5 & 2'h3 == row_5 ? 4'h2 : _GEN_202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_204 = 4'h3 == col_5 & 2'h0 == row_5 ? 4'hf : _GEN_203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_205 = 4'h3 == col_5 & 2'h1 == row_5 ? 4'h2 : _GEN_204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_206 = 4'h3 == col_5 & 2'h2 == row_5 ? 4'h5 : _GEN_205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_207 = 4'h3 == col_5 & 2'h3 == row_5 ? 4'hc : _GEN_206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_208 = 4'h4 == col_5 & 2'h0 == row_5 ? 4'h9 : _GEN_207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_209 = 4'h4 == col_5 & 2'h1 == row_5 ? 4'h7 : _GEN_208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_210 = 4'h4 == col_5 & 2'h2 == row_5 ? 4'h2 : _GEN_209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_211 = 4'h4 == col_5 & 2'h3 == row_5 ? 4'h9 : _GEN_210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_212 = 4'h5 == col_5 & 2'h0 == row_5 ? 4'h2 : _GEN_211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_213 = 4'h5 == col_5 & 2'h1 == row_5 ? 4'hc : _GEN_212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_214 = 4'h5 == col_5 & 2'h2 == row_5 ? 4'h8 : _GEN_213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_215 = 4'h5 == col_5 & 2'h3 == row_5 ? 4'h5 : _GEN_214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_216 = 4'h6 == col_5 & 2'h0 == row_5 ? 4'h6 : _GEN_215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_217 = 4'h6 == col_5 & 2'h1 == row_5 ? 4'h9 : _GEN_216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_218 = 4'h6 == col_5 & 2'h2 == row_5 ? 4'hc : _GEN_217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_219 = 4'h6 == col_5 & 2'h3 == row_5 ? 4'hf : _GEN_218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_220 = 4'h7 == col_5 & 2'h0 == row_5 ? 4'h8 : _GEN_219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_221 = 4'h7 == col_5 & 2'h1 == row_5 ? 4'h5 : _GEN_220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_222 = 4'h7 == col_5 & 2'h2 == row_5 ? 4'h3 : _GEN_221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_223 = 4'h7 == col_5 & 2'h3 == row_5 ? 4'ha : _GEN_222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_224 = 4'h8 == col_5 & 2'h0 == row_5 ? 4'h0 : _GEN_223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_225 = 4'h8 == col_5 & 2'h1 == row_5 ? 4'h6 : _GEN_224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_226 = 4'h8 == col_5 & 2'h2 == row_5 ? 4'h7 : _GEN_225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_227 = 4'h8 == col_5 & 2'h3 == row_5 ? 4'hb : _GEN_226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_228 = 4'h9 == col_5 & 2'h0 == row_5 ? 4'hd : _GEN_227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_229 = 4'h9 == col_5 & 2'h1 == row_5 ? 4'h1 : _GEN_228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_230 = 4'h9 == col_5 & 2'h2 == row_5 ? 4'h0 : _GEN_229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_231 = 4'h9 == col_5 & 2'h3 == row_5 ? 4'he : _GEN_230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_232 = 4'ha == col_5 & 2'h0 == row_5 ? 4'h3 : _GEN_231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_233 = 4'ha == col_5 & 2'h1 == row_5 ? 4'hd : _GEN_232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_234 = 4'ha == col_5 & 2'h2 == row_5 ? 4'h4 : _GEN_233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_235 = 4'ha == col_5 & 2'h3 == row_5 ? 4'h1 : _GEN_234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_236 = 4'hb == col_5 & 2'h0 == row_5 ? 4'h4 : _GEN_235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_237 = 4'hb == col_5 & 2'h1 == row_5 ? 4'he : _GEN_236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_238 = 4'hb == col_5 & 2'h2 == row_5 ? 4'ha : _GEN_237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_239 = 4'hb == col_5 & 2'h3 == row_5 ? 4'h7 : _GEN_238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_240 = 4'hc == col_5 & 2'h0 == row_5 ? 4'he : _GEN_239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_241 = 4'hc == col_5 & 2'h1 == row_5 ? 4'h0 : _GEN_240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_242 = 4'hc == col_5 & 2'h2 == row_5 ? 4'h1 : _GEN_241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_243 = 4'hc == col_5 & 2'h3 == row_5 ? 4'h6 : _GEN_242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_244 = 4'hd == col_5 & 2'h0 == row_5 ? 4'h7 : _GEN_243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_245 = 4'hd == col_5 & 2'h1 == row_5 ? 4'hb : _GEN_244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_246 = 4'hd == col_5 & 2'h2 == row_5 ? 4'hd : _GEN_245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_247 = 4'hd == col_5 & 2'h3 == row_5 ? 4'h0 : _GEN_246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_248 = 4'he == col_5 & 2'h0 == row_5 ? 4'h5 : _GEN_247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_249 = 4'he == col_5 & 2'h1 == row_5 ? 4'h3 : _GEN_248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_250 = 4'he == col_5 & 2'h2 == row_5 ? 4'hb : _GEN_249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_251 = 4'he == col_5 & 2'h3 == row_5 ? 4'h8 : _GEN_250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_252 = 4'hf == col_5 & 2'h0 == row_5 ? 4'hb : _GEN_251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_253 = 4'hf == col_5 & 2'h1 == row_5 ? 4'h8 : _GEN_252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_254 = 4'hf == col_5 & 2'h2 == row_5 ? 4'h6 : _GEN_253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_255 = 4'hf == col_5 & 2'h3 == row_5 ? 4'hd : _GEN_254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [15:0] lo_8 = {_GEN_191,_GEN_255,_GEN_63,_GEN_127}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_257 = 4'h0 == col_2 & 2'h1 == row_2 ? 4'hd : 4'ha; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_258 = 4'h0 == col_2 & 2'h2 == row_2 ? 4'hd : _GEN_257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_259 = 4'h0 == col_2 & 2'h3 == row_2 ? 4'h1 : _GEN_258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_260 = 4'h1 == col_2 & 2'h0 == row_2 ? 4'h0 : _GEN_259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_261 = 4'h1 == col_2 & 2'h1 == row_2 ? 4'h7 : _GEN_260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_262 = 4'h1 == col_2 & 2'h2 == row_2 ? 4'h6 : _GEN_261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_263 = 4'h1 == col_2 & 2'h3 == row_2 ? 4'ha : _GEN_262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_264 = 4'h2 == col_2 & 2'h0 == row_2 ? 4'h9 : _GEN_263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_265 = 4'h2 == col_2 & 2'h1 == row_2 ? 4'h0 : _GEN_264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_266 = 4'h2 == col_2 & 2'h2 == row_2 ? 4'h4 : _GEN_265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_267 = 4'h2 == col_2 & 2'h3 == row_2 ? 4'hd : _GEN_266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_268 = 4'h3 == col_2 & 2'h0 == row_2 ? 4'he : _GEN_267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_269 = 4'h3 == col_2 & 2'h1 == row_2 ? 4'h9 : _GEN_268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_270 = 4'h3 == col_2 & 2'h2 == row_2 ? 4'h9 : _GEN_269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_271 = 4'h3 == col_2 & 2'h3 == row_2 ? 4'h0 : _GEN_270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_272 = 4'h4 == col_2 & 2'h0 == row_2 ? 4'h6 : _GEN_271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_273 = 4'h4 == col_2 & 2'h1 == row_2 ? 4'h3 : _GEN_272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_274 = 4'h4 == col_2 & 2'h2 == row_2 ? 4'h8 : _GEN_273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_275 = 4'h4 == col_2 & 2'h3 == row_2 ? 4'h6 : _GEN_274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_276 = 4'h5 == col_2 & 2'h0 == row_2 ? 4'h3 : _GEN_275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_277 = 4'h5 == col_2 & 2'h1 == row_2 ? 4'h4 : _GEN_276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_278 = 4'h5 == col_2 & 2'h2 == row_2 ? 4'hf : _GEN_277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_279 = 4'h5 == col_2 & 2'h3 == row_2 ? 4'h9 : _GEN_278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_280 = 4'h6 == col_2 & 2'h0 == row_2 ? 4'hf : _GEN_279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_281 = 4'h6 == col_2 & 2'h1 == row_2 ? 4'h6 : _GEN_280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_282 = 4'h6 == col_2 & 2'h2 == row_2 ? 4'h3 : _GEN_281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_283 = 4'h6 == col_2 & 2'h3 == row_2 ? 4'h8 : _GEN_282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_284 = 4'h7 == col_2 & 2'h0 == row_2 ? 4'h5 : _GEN_283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_285 = 4'h7 == col_2 & 2'h1 == row_2 ? 4'ha : _GEN_284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_286 = 4'h7 == col_2 & 2'h2 == row_2 ? 4'h0 : _GEN_285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_287 = 4'h7 == col_2 & 2'h3 == row_2 ? 4'h7 : _GEN_286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_288 = 4'h8 == col_2 & 2'h0 == row_2 ? 4'h1 : _GEN_287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_289 = 4'h8 == col_2 & 2'h1 == row_2 ? 4'h2 : _GEN_288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_290 = 4'h8 == col_2 & 2'h2 == row_2 ? 4'hb : _GEN_289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_291 = 4'h8 == col_2 & 2'h3 == row_2 ? 4'h4 : _GEN_290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_292 = 4'h9 == col_2 & 2'h0 == row_2 ? 4'hd : _GEN_291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_293 = 4'h9 == col_2 & 2'h1 == row_2 ? 4'h8 : _GEN_292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_294 = 4'h9 == col_2 & 2'h2 == row_2 ? 4'h1 : _GEN_293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_295 = 4'h9 == col_2 & 2'h3 == row_2 ? 4'hf : _GEN_294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_296 = 4'ha == col_2 & 2'h0 == row_2 ? 4'hc : _GEN_295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_297 = 4'ha == col_2 & 2'h1 == row_2 ? 4'h5 : _GEN_296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_298 = 4'ha == col_2 & 2'h2 == row_2 ? 4'h2 : _GEN_297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_299 = 4'ha == col_2 & 2'h3 == row_2 ? 4'he : _GEN_298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_300 = 4'hb == col_2 & 2'h0 == row_2 ? 4'h7 : _GEN_299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_301 = 4'hb == col_2 & 2'h1 == row_2 ? 4'he : _GEN_300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_302 = 4'hb == col_2 & 2'h2 == row_2 ? 4'hc : _GEN_301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_303 = 4'hb == col_2 & 2'h3 == row_2 ? 4'h3 : _GEN_302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_304 = 4'hc == col_2 & 2'h0 == row_2 ? 4'hb : _GEN_303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_305 = 4'hc == col_2 & 2'h1 == row_2 ? 4'hc : _GEN_304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_306 = 4'hc == col_2 & 2'h2 == row_2 ? 4'h5 : _GEN_305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_307 = 4'hc == col_2 & 2'h3 == row_2 ? 4'hb : _GEN_306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_308 = 4'hd == col_2 & 2'h0 == row_2 ? 4'h4 : _GEN_307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_309 = 4'hd == col_2 & 2'h1 == row_2 ? 4'hb : _GEN_308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_310 = 4'hd == col_2 & 2'h2 == row_2 ? 4'ha : _GEN_309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_311 = 4'hd == col_2 & 2'h3 == row_2 ? 4'h5 : _GEN_310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_312 = 4'he == col_2 & 2'h0 == row_2 ? 4'h2 : _GEN_311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_313 = 4'he == col_2 & 2'h1 == row_2 ? 4'hf : _GEN_312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_314 = 4'he == col_2 & 2'h2 == row_2 ? 4'he : _GEN_313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_315 = 4'he == col_2 & 2'h3 == row_2 ? 4'h2 : _GEN_314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_316 = 4'hf == col_2 & 2'h0 == row_2 ? 4'h8 : _GEN_315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_317 = 4'hf == col_2 & 2'h1 == row_2 ? 4'h1 : _GEN_316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_318 = 4'hf == col_2 & 2'h2 == row_2 ? 4'h7 : _GEN_317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_319 = 4'hf == col_2 & 2'h3 == row_2 ? 4'hc : _GEN_318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_321 = 4'h0 == col_3 & 2'h1 == row_3 ? 4'hd : 4'h7; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_322 = 4'h0 == col_3 & 2'h2 == row_3 ? 4'ha : _GEN_321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_323 = 4'h0 == col_3 & 2'h3 == row_3 ? 4'h3 : _GEN_322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_324 = 4'h1 == col_3 & 2'h0 == row_3 ? 4'hd : _GEN_323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_325 = 4'h1 == col_3 & 2'h1 == row_3 ? 4'h8 : _GEN_324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_326 = 4'h1 == col_3 & 2'h2 == row_3 ? 4'h6 : _GEN_325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_327 = 4'h1 == col_3 & 2'h3 == row_3 ? 4'hf : _GEN_326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_328 = 4'h2 == col_3 & 2'h0 == row_3 ? 4'he : _GEN_327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_329 = 4'h2 == col_3 & 2'h1 == row_3 ? 4'hb : _GEN_328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_330 = 4'h2 == col_3 & 2'h2 == row_3 ? 4'h9 : _GEN_329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_331 = 4'h2 == col_3 & 2'h3 == row_3 ? 4'h0 : _GEN_330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_332 = 4'h3 == col_3 & 2'h0 == row_3 ? 4'h3 : _GEN_331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_333 = 4'h3 == col_3 & 2'h1 == row_3 ? 4'h5 : _GEN_332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_334 = 4'h3 == col_3 & 2'h2 == row_3 ? 4'h0 : _GEN_333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_335 = 4'h3 == col_3 & 2'h3 == row_3 ? 4'h6 : _GEN_334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_336 = 4'h4 == col_3 & 2'h0 == row_3 ? 4'h0 : _GEN_335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_337 = 4'h4 == col_3 & 2'h1 == row_3 ? 4'h6 : _GEN_336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_338 = 4'h4 == col_3 & 2'h2 == row_3 ? 4'hc : _GEN_337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_339 = 4'h4 == col_3 & 2'h3 == row_3 ? 4'ha : _GEN_338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_340 = 4'h5 == col_3 & 2'h0 == row_3 ? 4'h6 : _GEN_339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_341 = 4'h5 == col_3 & 2'h1 == row_3 ? 4'hf : _GEN_340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_342 = 4'h5 == col_3 & 2'h2 == row_3 ? 4'hb : _GEN_341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_343 = 4'h5 == col_3 & 2'h3 == row_3 ? 4'h1 : _GEN_342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_344 = 4'h6 == col_3 & 2'h0 == row_3 ? 4'h9 : _GEN_343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_345 = 4'h6 == col_3 & 2'h1 == row_3 ? 4'h0 : _GEN_344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_346 = 4'h6 == col_3 & 2'h2 == row_3 ? 4'h7 : _GEN_345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_347 = 4'h6 == col_3 & 2'h3 == row_3 ? 4'hd : _GEN_346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_348 = 4'h7 == col_3 & 2'h0 == row_3 ? 4'ha : _GEN_347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_349 = 4'h7 == col_3 & 2'h1 == row_3 ? 4'h3 : _GEN_348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_350 = 4'h7 == col_3 & 2'h2 == row_3 ? 4'hd : _GEN_349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_351 = 4'h7 == col_3 & 2'h3 == row_3 ? 4'h8 : _GEN_350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_352 = 4'h8 == col_3 & 2'h0 == row_3 ? 4'h1 : _GEN_351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_353 = 4'h8 == col_3 & 2'h1 == row_3 ? 4'h4 : _GEN_352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_354 = 4'h8 == col_3 & 2'h2 == row_3 ? 4'hf : _GEN_353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_355 = 4'h8 == col_3 & 2'h3 == row_3 ? 4'h9 : _GEN_354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_356 = 4'h9 == col_3 & 2'h0 == row_3 ? 4'h2 : _GEN_355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_357 = 4'h9 == col_3 & 2'h1 == row_3 ? 4'h7 : _GEN_356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_358 = 4'h9 == col_3 & 2'h2 == row_3 ? 4'h1 : _GEN_357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_359 = 4'h9 == col_3 & 2'h3 == row_3 ? 4'h4 : _GEN_358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_360 = 4'ha == col_3 & 2'h0 == row_3 ? 4'h8 : _GEN_359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_361 = 4'ha == col_3 & 2'h1 == row_3 ? 4'h2 : _GEN_360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_362 = 4'ha == col_3 & 2'h2 == row_3 ? 4'h3 : _GEN_361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_363 = 4'ha == col_3 & 2'h3 == row_3 ? 4'h5 : _GEN_362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_364 = 4'hb == col_3 & 2'h0 == row_3 ? 4'h5 : _GEN_363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_365 = 4'hb == col_3 & 2'h1 == row_3 ? 4'hc : _GEN_364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_366 = 4'hb == col_3 & 2'h2 == row_3 ? 4'he : _GEN_365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_367 = 4'hb == col_3 & 2'h3 == row_3 ? 4'hb : _GEN_366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_368 = 4'hc == col_3 & 2'h0 == row_3 ? 4'hb : _GEN_367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_369 = 4'hc == col_3 & 2'h1 == row_3 ? 4'h1 : _GEN_368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_370 = 4'hc == col_3 & 2'h2 == row_3 ? 4'h5 : _GEN_369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_371 = 4'hc == col_3 & 2'h3 == row_3 ? 4'hc : _GEN_370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_372 = 4'hd == col_3 & 2'h0 == row_3 ? 4'hc : _GEN_371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_373 = 4'hd == col_3 & 2'h1 == row_3 ? 4'ha : _GEN_372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_374 = 4'hd == col_3 & 2'h2 == row_3 ? 4'h2 : _GEN_373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_375 = 4'hd == col_3 & 2'h3 == row_3 ? 4'h7 : _GEN_374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_376 = 4'he == col_3 & 2'h0 == row_3 ? 4'h4 : _GEN_375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_377 = 4'he == col_3 & 2'h1 == row_3 ? 4'he : _GEN_376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_378 = 4'he == col_3 & 2'h2 == row_3 ? 4'h8 : _GEN_377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_379 = 4'he == col_3 & 2'h3 == row_3 ? 4'h2 : _GEN_378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_380 = 4'hf == col_3 & 2'h0 == row_3 ? 4'hf : _GEN_379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_381 = 4'hf == col_3 & 2'h1 == row_3 ? 4'h9 : _GEN_380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_382 = 4'hf == col_3 & 2'h2 == row_3 ? 4'h4 : _GEN_381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_383 = 4'hf == col_3 & 2'h3 == row_3 ? 4'he : _GEN_382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_385 = 4'h0 == col_0 & 2'h1 == row_0 ? 4'h0 : 4'he; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_386 = 4'h0 == col_0 & 2'h2 == row_0 ? 4'h4 : _GEN_385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_387 = 4'h0 == col_0 & 2'h3 == row_0 ? 4'hf : _GEN_386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_388 = 4'h1 == col_0 & 2'h0 == row_0 ? 4'h4 : _GEN_387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_389 = 4'h1 == col_0 & 2'h1 == row_0 ? 4'hf : _GEN_388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_390 = 4'h1 == col_0 & 2'h2 == row_0 ? 4'h1 : _GEN_389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_391 = 4'h1 == col_0 & 2'h3 == row_0 ? 4'hc : _GEN_390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_392 = 4'h2 == col_0 & 2'h0 == row_0 ? 4'hd : _GEN_391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_393 = 4'h2 == col_0 & 2'h1 == row_0 ? 4'h7 : _GEN_392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_394 = 4'h2 == col_0 & 2'h2 == row_0 ? 4'he : _GEN_393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_395 = 4'h2 == col_0 & 2'h3 == row_0 ? 4'h8 : _GEN_394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_396 = 4'h3 == col_0 & 2'h0 == row_0 ? 4'h1 : _GEN_395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_397 = 4'h3 == col_0 & 2'h1 == row_0 ? 4'h4 : _GEN_396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_398 = 4'h3 == col_0 & 2'h2 == row_0 ? 4'h8 : _GEN_397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_399 = 4'h3 == col_0 & 2'h3 == row_0 ? 4'h2 : _GEN_398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_400 = 4'h4 == col_0 & 2'h0 == row_0 ? 4'h2 : _GEN_399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_401 = 4'h4 == col_0 & 2'h1 == row_0 ? 4'he : _GEN_400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_402 = 4'h4 == col_0 & 2'h2 == row_0 ? 4'hd : _GEN_401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_403 = 4'h4 == col_0 & 2'h3 == row_0 ? 4'h4 : _GEN_402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_404 = 4'h5 == col_0 & 2'h0 == row_0 ? 4'hf : _GEN_403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_405 = 4'h5 == col_0 & 2'h1 == row_0 ? 4'h2 : _GEN_404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_406 = 4'h5 == col_0 & 2'h2 == row_0 ? 4'h6 : _GEN_405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_407 = 4'h5 == col_0 & 2'h3 == row_0 ? 4'h9 : _GEN_406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_408 = 4'h6 == col_0 & 2'h0 == row_0 ? 4'hb : _GEN_407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_409 = 4'h6 == col_0 & 2'h1 == row_0 ? 4'hd : _GEN_408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_410 = 4'h6 == col_0 & 2'h2 == row_0 ? 4'h2 : _GEN_409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_411 = 4'h6 == col_0 & 2'h3 == row_0 ? 4'h1 : _GEN_410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_412 = 4'h7 == col_0 & 2'h0 == row_0 ? 4'h8 : _GEN_411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_413 = 4'h7 == col_0 & 2'h1 == row_0 ? 4'h1 : _GEN_412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_414 = 4'h7 == col_0 & 2'h2 == row_0 ? 4'hb : _GEN_413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_415 = 4'h7 == col_0 & 2'h3 == row_0 ? 4'h7 : _GEN_414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_416 = 4'h8 == col_0 & 2'h0 == row_0 ? 4'h3 : _GEN_415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_417 = 4'h8 == col_0 & 2'h1 == row_0 ? 4'ha : _GEN_416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_418 = 4'h8 == col_0 & 2'h2 == row_0 ? 4'hf : _GEN_417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_419 = 4'h8 == col_0 & 2'h3 == row_0 ? 4'h5 : _GEN_418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_420 = 4'h9 == col_0 & 2'h0 == row_0 ? 4'ha : _GEN_419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_421 = 4'h9 == col_0 & 2'h1 == row_0 ? 4'h6 : _GEN_420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_422 = 4'h9 == col_0 & 2'h2 == row_0 ? 4'hc : _GEN_421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_423 = 4'h9 == col_0 & 2'h3 == row_0 ? 4'hb : _GEN_422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_424 = 4'ha == col_0 & 2'h0 == row_0 ? 4'h6 : _GEN_423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_425 = 4'ha == col_0 & 2'h1 == row_0 ? 4'hc : _GEN_424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_426 = 4'ha == col_0 & 2'h2 == row_0 ? 4'h9 : _GEN_425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_427 = 4'ha == col_0 & 2'h3 == row_0 ? 4'h3 : _GEN_426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_428 = 4'hb == col_0 & 2'h0 == row_0 ? 4'hc : _GEN_427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_429 = 4'hb == col_0 & 2'h1 == row_0 ? 4'hb : _GEN_428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_430 = 4'hb == col_0 & 2'h2 == row_0 ? 4'h7 : _GEN_429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_431 = 4'hb == col_0 & 2'h3 == row_0 ? 4'he : _GEN_430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_432 = 4'hc == col_0 & 2'h0 == row_0 ? 4'h5 : _GEN_431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_433 = 4'hc == col_0 & 2'h1 == row_0 ? 4'h9 : _GEN_432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_434 = 4'hc == col_0 & 2'h2 == row_0 ? 4'h3 : _GEN_433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_435 = 4'hc == col_0 & 2'h3 == row_0 ? 4'ha : _GEN_434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_436 = 4'hd == col_0 & 2'h0 == row_0 ? 4'h9 : _GEN_435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_437 = 4'hd == col_0 & 2'h1 == row_0 ? 4'h5 : _GEN_436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_438 = 4'hd == col_0 & 2'h2 == row_0 ? 4'ha : _GEN_437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_439 = 4'hd == col_0 & 2'h3 == row_0 ? 4'h0 : _GEN_438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_440 = 4'he == col_0 & 2'h0 == row_0 ? 4'h0 : _GEN_439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_441 = 4'he == col_0 & 2'h1 == row_0 ? 4'h3 : _GEN_440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_442 = 4'he == col_0 & 2'h2 == row_0 ? 4'h5 : _GEN_441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_443 = 4'he == col_0 & 2'h3 == row_0 ? 4'h6 : _GEN_442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_444 = 4'hf == col_0 & 2'h0 == row_0 ? 4'h7 : _GEN_443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_445 = 4'hf == col_0 & 2'h1 == row_0 ? 4'h8 : _GEN_444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_446 = 4'hf == col_0 & 2'h2 == row_0 ? 4'h0 : _GEN_445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_447 = 4'hf == col_0 & 2'h3 == row_0 ? 4'hd : _GEN_446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_449 = 4'h0 == col_1 & 2'h1 == row_1 ? 4'h3 : 4'hf; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_450 = 4'h0 == col_1 & 2'h2 == row_1 ? 4'h0 : _GEN_449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_451 = 4'h0 == col_1 & 2'h3 == row_1 ? 4'hd : _GEN_450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_452 = 4'h1 == col_1 & 2'h0 == row_1 ? 4'h1 : _GEN_451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_453 = 4'h1 == col_1 & 2'h1 == row_1 ? 4'hd : _GEN_452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_454 = 4'h1 == col_1 & 2'h2 == row_1 ? 4'he : _GEN_453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_455 = 4'h1 == col_1 & 2'h3 == row_1 ? 4'h8 : _GEN_454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_456 = 4'h2 == col_1 & 2'h0 == row_1 ? 4'h8 : _GEN_455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_457 = 4'h2 == col_1 & 2'h1 == row_1 ? 4'h4 : _GEN_456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_458 = 4'h2 == col_1 & 2'h2 == row_1 ? 4'h7 : _GEN_457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_459 = 4'h2 == col_1 & 2'h3 == row_1 ? 4'ha : _GEN_458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_460 = 4'h3 == col_1 & 2'h0 == row_1 ? 4'he : _GEN_459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_461 = 4'h3 == col_1 & 2'h1 == row_1 ? 4'h7 : _GEN_460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_462 = 4'h3 == col_1 & 2'h2 == row_1 ? 4'hb : _GEN_461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_463 = 4'h3 == col_1 & 2'h3 == row_1 ? 4'h1 : _GEN_462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_464 = 4'h4 == col_1 & 2'h0 == row_1 ? 4'h6 : _GEN_463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_465 = 4'h4 == col_1 & 2'h1 == row_1 ? 4'hf : _GEN_464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_466 = 4'h4 == col_1 & 2'h2 == row_1 ? 4'ha : _GEN_465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_467 = 4'h4 == col_1 & 2'h3 == row_1 ? 4'h3 : _GEN_466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_468 = 4'h5 == col_1 & 2'h0 == row_1 ? 4'hb : _GEN_467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_469 = 4'h5 == col_1 & 2'h1 == row_1 ? 4'h2 : _GEN_468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_470 = 4'h5 == col_1 & 2'h2 == row_1 ? 4'h4 : _GEN_469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_471 = 4'h5 == col_1 & 2'h3 == row_1 ? 4'hf : _GEN_470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_472 = 4'h6 == col_1 & 2'h0 == row_1 ? 4'h3 : _GEN_471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_473 = 4'h6 == col_1 & 2'h1 == row_1 ? 4'h8 : _GEN_472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_474 = 4'h6 == col_1 & 2'h2 == row_1 ? 4'hd : _GEN_473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_475 = 4'h6 == col_1 & 2'h3 == row_1 ? 4'h4 : _GEN_474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_476 = 4'h7 == col_1 & 2'h0 == row_1 ? 4'h4 : _GEN_475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_477 = 4'h7 == col_1 & 2'h1 == row_1 ? 4'he : _GEN_476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_478 = 4'h7 == col_1 & 2'h2 == row_1 ? 4'h1 : _GEN_477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_479 = 4'h7 == col_1 & 2'h3 == row_1 ? 4'h2 : _GEN_478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_480 = 4'h8 == col_1 & 2'h0 == row_1 ? 4'h9 : _GEN_479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_481 = 4'h8 == col_1 & 2'h1 == row_1 ? 4'hc : _GEN_480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_482 = 4'h8 == col_1 & 2'h2 == row_1 ? 4'h5 : _GEN_481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_483 = 4'h8 == col_1 & 2'h3 == row_1 ? 4'hb : _GEN_482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_484 = 4'h9 == col_1 & 2'h0 == row_1 ? 4'h7 : _GEN_483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_485 = 4'h9 == col_1 & 2'h1 == row_1 ? 4'h0 : _GEN_484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_486 = 4'h9 == col_1 & 2'h2 == row_1 ? 4'h8 : _GEN_485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_487 = 4'h9 == col_1 & 2'h3 == row_1 ? 4'h6 : _GEN_486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_488 = 4'ha == col_1 & 2'h0 == row_1 ? 4'h2 : _GEN_487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_489 = 4'ha == col_1 & 2'h1 == row_1 ? 4'h1 : _GEN_488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_490 = 4'ha == col_1 & 2'h2 == row_1 ? 4'hc : _GEN_489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_491 = 4'ha == col_1 & 2'h3 == row_1 ? 4'h7 : _GEN_490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_492 = 4'hb == col_1 & 2'h0 == row_1 ? 4'hd : _GEN_491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_493 = 4'hb == col_1 & 2'h1 == row_1 ? 4'ha : _GEN_492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_494 = 4'hb == col_1 & 2'h2 == row_1 ? 4'h6 : _GEN_493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_495 = 4'hb == col_1 & 2'h3 == row_1 ? 4'hc : _GEN_494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_496 = 4'hc == col_1 & 2'h0 == row_1 ? 4'hc : _GEN_495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_497 = 4'hc == col_1 & 2'h1 == row_1 ? 4'h6 : _GEN_496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_498 = 4'hc == col_1 & 2'h2 == row_1 ? 4'h9 : _GEN_497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_499 = 4'hc == col_1 & 2'h3 == row_1 ? 4'h0 : _GEN_498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_500 = 4'hd == col_1 & 2'h0 == row_1 ? 4'h0 : _GEN_499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_501 = 4'hd == col_1 & 2'h1 == row_1 ? 4'h9 : _GEN_500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_502 = 4'hd == col_1 & 2'h2 == row_1 ? 4'h3 : _GEN_501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_503 = 4'hd == col_1 & 2'h3 == row_1 ? 4'h5 : _GEN_502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_504 = 4'he == col_1 & 2'h0 == row_1 ? 4'h5 : _GEN_503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_505 = 4'he == col_1 & 2'h1 == row_1 ? 4'hb : _GEN_504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_506 = 4'he == col_1 & 2'h2 == row_1 ? 4'h2 : _GEN_505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_507 = 4'he == col_1 & 2'h3 == row_1 ? 4'he : _GEN_506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_508 = 4'hf == col_1 & 2'h0 == row_1 ? 4'ha : _GEN_507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_509 = 4'hf == col_1 & 2'h1 == row_1 ? 4'h5 : _GEN_508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_510 = 4'hf == col_1 & 2'h2 == row_1 ? 4'hf : _GEN_509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [3:0] _GEN_511 = 4'hf == col_1 & 2'h3 == row_1 ? 4'h9 : _GEN_510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [15:0] hi_8 = {_GEN_447,_GEN_511,_GEN_319,_GEN_383}; // @[Cat.scala 30:58]
  assign io_out = {hi_8,lo_8}; // @[Cat.scala 30:58]
endmodule
module DES_P(
  input  [31:0] io_in,
  output [31:0] io_out
);
  wire [31:0] _T_3 = {{16'd0}, io_in[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_5 = {io_in[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_7 = _T_5 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_8 = _T_3 | _T_7; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_0 = {{8'd0}, _T_8[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_13 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_15 = {_T_8[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_17 = _T_15 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_18 = _T_13 | _T_17; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1 = {{4'd0}, _T_18[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_23 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_25 = {_T_18[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_27 = _T_25 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_28 = _T_23 | _T_27; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_2 = {{2'd0}, _T_28[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_33 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_35 = {_T_28[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_37 = _T_35 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_38 = _T_33 | _T_37; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3 = {{1'd0}, _T_38[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_43 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_45 = {_T_38[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_47 = _T_45 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] reversed = _T_43 | _T_47; // @[Bitwise.scala 103:39]
  wire  hi_hi_hi_hi_hi = reversed[15]; // @[DES_FSM.scala 475:25]
  wire  hi_hi_hi_hi_lo = reversed[6]; // @[DES_FSM.scala 475:38]
  wire  hi_hi_hi_lo_hi = reversed[19]; // @[DES_FSM.scala 475:50]
  wire  hi_hi_hi_lo_lo = reversed[20]; // @[DES_FSM.scala 475:63]
  wire  hi_hi_lo_hi_hi = reversed[28]; // @[DES_FSM.scala 476:13]
  wire  hi_hi_lo_hi_lo = reversed[11]; // @[DES_FSM.scala 476:26]
  wire  hi_hi_lo_lo_hi = reversed[27]; // @[DES_FSM.scala 476:39]
  wire  hi_hi_lo_lo_lo = reversed[16]; // @[DES_FSM.scala 476:52]
  wire  hi_lo_hi_hi_hi = reversed[0]; // @[DES_FSM.scala 477:13]
  wire  hi_lo_hi_hi_lo = reversed[14]; // @[DES_FSM.scala 477:25]
  wire  hi_lo_hi_lo_hi = reversed[22]; // @[DES_FSM.scala 477:38]
  wire  hi_lo_hi_lo_lo = reversed[25]; // @[DES_FSM.scala 477:51]
  wire  hi_lo_lo_hi_hi = reversed[4]; // @[DES_FSM.scala 478:13]
  wire  hi_lo_lo_hi_lo = reversed[17]; // @[DES_FSM.scala 478:25]
  wire  hi_lo_lo_lo_hi = reversed[30]; // @[DES_FSM.scala 478:38]
  wire  hi_lo_lo_lo_lo = reversed[9]; // @[DES_FSM.scala 478:51]
  wire  lo_hi_hi_hi_hi = reversed[1]; // @[DES_FSM.scala 479:13]
  wire  lo_hi_hi_hi_lo = reversed[7]; // @[DES_FSM.scala 479:25]
  wire  lo_hi_hi_lo_hi = reversed[23]; // @[DES_FSM.scala 479:37]
  wire  lo_hi_hi_lo_lo = reversed[13]; // @[DES_FSM.scala 479:50]
  wire  lo_hi_lo_hi_hi = reversed[31]; // @[DES_FSM.scala 480:13]
  wire  lo_hi_lo_hi_lo = reversed[26]; // @[DES_FSM.scala 480:26]
  wire  lo_hi_lo_lo_hi = reversed[2]; // @[DES_FSM.scala 480:39]
  wire  lo_hi_lo_lo_lo = reversed[8]; // @[DES_FSM.scala 480:51]
  wire  lo_lo_hi_hi_hi = reversed[18]; // @[DES_FSM.scala 481:13]
  wire  lo_lo_hi_hi_lo = reversed[12]; // @[DES_FSM.scala 481:26]
  wire  lo_lo_hi_lo_hi = reversed[29]; // @[DES_FSM.scala 481:39]
  wire  lo_lo_hi_lo_lo = reversed[5]; // @[DES_FSM.scala 481:52]
  wire  lo_lo_lo_hi_hi = reversed[21]; // @[DES_FSM.scala 482:13]
  wire  lo_lo_lo_hi_lo = reversed[10]; // @[DES_FSM.scala 482:26]
  wire  lo_lo_lo_lo_hi = reversed[3]; // @[DES_FSM.scala 482:39]
  wire  lo_lo_lo_lo_lo = reversed[24]; // @[DES_FSM.scala 482:51]
  wire [7:0] lo_lo = {lo_lo_hi_hi_hi,lo_lo_hi_hi_lo,lo_lo_hi_lo_hi,lo_lo_hi_lo_lo,lo_lo_lo_hi_hi,lo_lo_lo_hi_lo,
    lo_lo_lo_lo_hi,lo_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [15:0] lo = {lo_hi_hi_hi_hi,lo_hi_hi_hi_lo,lo_hi_hi_lo_hi,lo_hi_hi_lo_lo,lo_hi_lo_hi_hi,lo_hi_lo_hi_lo,
    lo_hi_lo_lo_hi,lo_hi_lo_lo_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo = {hi_lo_hi_hi_hi,hi_lo_hi_hi_lo,hi_lo_hi_lo_hi,hi_lo_hi_lo_lo,hi_lo_lo_hi_hi,hi_lo_lo_hi_lo,
    hi_lo_lo_lo_hi,hi_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [15:0] hi = {hi_hi_hi_hi_hi,hi_hi_hi_hi_lo,hi_hi_hi_lo_hi,hi_hi_hi_lo_lo,hi_hi_lo_hi_hi,hi_hi_lo_hi_lo,
    hi_hi_lo_lo_hi,hi_hi_lo_lo_lo,hi_lo}; // @[Cat.scala 30:58]
  assign io_out = {hi,lo}; // @[Cat.scala 30:58]
endmodule
module DES_f(
  input  [31:0] io_R,
  input  [47:0] io_K,
  output [31:0] io_out
);
  wire [31:0] E_io_R; // @[DES_FSM.scala 300:17]
  wire [47:0] E_io_E; // @[DES_FSM.scala 300:17]
  wire [47:0] S_io_in; // @[DES_FSM.scala 303:17]
  wire [31:0] S_io_out; // @[DES_FSM.scala 303:17]
  wire [31:0] P_io_in; // @[DES_FSM.scala 306:17]
  wire [31:0] P_io_out; // @[DES_FSM.scala 306:17]
  DES_E E ( // @[DES_FSM.scala 300:17]
    .io_R(E_io_R),
    .io_E(E_io_E)
  );
  DES_S S ( // @[DES_FSM.scala 303:17]
    .io_in(S_io_in),
    .io_out(S_io_out)
  );
  DES_P P ( // @[DES_FSM.scala 306:17]
    .io_in(P_io_in),
    .io_out(P_io_out)
  );
  assign io_out = P_io_out; // @[DES_FSM.scala 308:10]
  assign E_io_R = io_R; // @[DES_FSM.scala 301:10]
  assign S_io_in = E_io_E ^ io_K; // @[DES_FSM.scala 304:21]
  assign P_io_in = S_io_out; // @[DES_FSM.scala 307:11]
endmodule
module DES_ProcessingElement(
  input  [4:0]  io_round,
  input  [31:0] io_in_L,
  input  [31:0] io_in_R,
  input  [27:0] io_in_C,
  input  [27:0] io_in_D,
  output [31:0] io_out_L,
  output [31:0] io_out_R,
  output [27:0] io_out_C,
  output [27:0] io_out_D
);
  wire [4:0] keys_io_round; // @[DES_FSM.scala 101:20]
  wire [27:0] keys_io_C; // @[DES_FSM.scala 101:20]
  wire [27:0] keys_io_D; // @[DES_FSM.scala 101:20]
  wire [27:0] keys_io_C_next; // @[DES_FSM.scala 101:20]
  wire [27:0] keys_io_D_next; // @[DES_FSM.scala 101:20]
  wire [47:0] keys_io_K; // @[DES_FSM.scala 101:20]
  wire [31:0] f_io_R; // @[DES_FSM.scala 106:17]
  wire [47:0] f_io_K; // @[DES_FSM.scala 106:17]
  wire [31:0] f_io_out; // @[DES_FSM.scala 106:17]
  DES_keys keys ( // @[DES_FSM.scala 101:20]
    .io_round(keys_io_round),
    .io_C(keys_io_C),
    .io_D(keys_io_D),
    .io_C_next(keys_io_C_next),
    .io_D_next(keys_io_D_next),
    .io_K(keys_io_K)
  );
  DES_f f ( // @[DES_FSM.scala 106:17]
    .io_R(f_io_R),
    .io_K(f_io_K),
    .io_out(f_io_out)
  );
  assign io_out_L = io_in_R; // @[DES_FSM.scala 110:12]
  assign io_out_R = io_in_L ^ f_io_out; // @[DES_FSM.scala 111:23]
  assign io_out_C = keys_io_C_next; // @[DES_FSM.scala 112:12]
  assign io_out_D = keys_io_D_next; // @[DES_FSM.scala 113:12]
  assign keys_io_round = io_round; // @[DES_FSM.scala 102:17]
  assign keys_io_C = io_in_C; // @[DES_FSM.scala 103:13]
  assign keys_io_D = io_in_D; // @[DES_FSM.scala 104:13]
  assign f_io_R = io_in_R; // @[DES_FSM.scala 107:10]
  assign f_io_K = keys_io_K; // @[DES_FSM.scala 108:10]
endmodule
module DES_FSM(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_text,
  input  [63:0] io_in_bits_key,
  input         io_result_ready,
  output        io_result_valid,
  output [63:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] ip_io_text; // @[DES_FSM.scala 27:18]
  wire [63:0] ip_io_key; // @[DES_FSM.scala 27:18]
  wire [31:0] ip_io_out_L; // @[DES_FSM.scala 27:18]
  wire [31:0] ip_io_out_R; // @[DES_FSM.scala 27:18]
  wire [27:0] ip_io_out_C; // @[DES_FSM.scala 27:18]
  wire [27:0] ip_io_out_D; // @[DES_FSM.scala 27:18]
  wire [31:0] fp_io_L; // @[DES_FSM.scala 30:18]
  wire [31:0] fp_io_R; // @[DES_FSM.scala 30:18]
  wire [63:0] fp_io_out; // @[DES_FSM.scala 30:18]
  wire [4:0] pe_io_round; // @[DES_FSM.scala 33:18]
  wire [31:0] pe_io_in_L; // @[DES_FSM.scala 33:18]
  wire [31:0] pe_io_in_R; // @[DES_FSM.scala 33:18]
  wire [27:0] pe_io_in_C; // @[DES_FSM.scala 33:18]
  wire [27:0] pe_io_in_D; // @[DES_FSM.scala 33:18]
  wire [31:0] pe_io_out_L; // @[DES_FSM.scala 33:18]
  wire [31:0] pe_io_out_R; // @[DES_FSM.scala 33:18]
  wire [27:0] pe_io_out_C; // @[DES_FSM.scala 33:18]
  wire [27:0] pe_io_out_D; // @[DES_FSM.scala 33:18]
  reg [2:0] stateReg; // @[DES_FSM.scala 16:25]
  reg [3:0] roundReg; // @[DES_FSM.scala 17:25]
  reg [63:0] textReg; // @[DES_FSM.scala 18:24]
  reg [63:0] keyReg; // @[DES_FSM.scala 19:23]
  reg [31:0] dataReg_L; // @[DES_FSM.scala 20:24]
  reg [31:0] dataReg_R; // @[DES_FSM.scala 20:24]
  reg [27:0] dataReg_C; // @[DES_FSM.scala 20:24]
  reg [27:0] dataReg_D; // @[DES_FSM.scala 20:24]
  reg [63:0] resultsReg; // @[DES_FSM.scala 21:27]
  wire  _T_2 = 3'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h2 == stateReg; // @[Conditional.scala 37:30]
  wire [3:0] _T_6 = roundReg + 4'h1; // @[DES_FSM.scala 55:28]
  wire [2:0] _GEN_3 = roundReg == 4'hf ? 3'h3 : stateReg; // @[DES_FSM.scala 56:31 DES_FSM.scala 57:18 DES_FSM.scala 16:25]
  wire  _T_8 = 3'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h4 == stateReg; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_4 = io_result_ready ? 3'h0 : stateReg; // @[DES_FSM.scala 67:29 DES_FSM.scala 68:18 DES_FSM.scala 16:25]
  wire [2:0] _GEN_5 = _T_9 ? _GEN_4 : stateReg; // @[Conditional.scala 39:67 DES_FSM.scala 16:25]
  wire [63:0] _GEN_8 = _T_8 ? fp_io_out : resultsReg; // @[Conditional.scala 39:67 DES_FSM.scala 63:18 DES_FSM.scala 21:27]
  wire [2:0] _GEN_9 = _T_8 ? 3'h4 : _GEN_5; // @[Conditional.scala 39:67 DES_FSM.scala 64:16]
  DES_InitialPermutation ip ( // @[DES_FSM.scala 27:18]
    .io_text(ip_io_text),
    .io_key(ip_io_key),
    .io_out_L(ip_io_out_L),
    .io_out_R(ip_io_out_R),
    .io_out_C(ip_io_out_C),
    .io_out_D(ip_io_out_D)
  );
  DES_FinalPermutation fp ( // @[DES_FSM.scala 30:18]
    .io_L(fp_io_L),
    .io_R(fp_io_R),
    .io_out(fp_io_out)
  );
  DES_ProcessingElement pe ( // @[DES_FSM.scala 33:18]
    .io_round(pe_io_round),
    .io_in_L(pe_io_in_L),
    .io_in_R(pe_io_in_R),
    .io_in_C(pe_io_in_C),
    .io_in_D(pe_io_in_D),
    .io_out_L(pe_io_out_L),
    .io_out_R(pe_io_out_R),
    .io_out_C(pe_io_out_C),
    .io_out_D(pe_io_out_D)
  );
  assign io_in_ready = stateReg == 3'h0; // @[DES_FSM.scala 23:27]
  assign io_result_valid = stateReg == 3'h4; // @[DES_FSM.scala 24:31]
  assign io_result_bits = resultsReg; // @[DES_FSM.scala 25:18]
  assign ip_io_text = textReg; // @[Conditional.scala 39:67 DES_FSM.scala 45:18]
  assign ip_io_key = keyReg; // @[Conditional.scala 39:67 DES_FSM.scala 46:17]
  assign fp_io_L = dataReg_L; // @[Conditional.scala 39:67 DES_FSM.scala 62:15]
  assign fp_io_R = dataReg_R; // @[Conditional.scala 39:67 DES_FSM.scala 61:15]
  assign pe_io_round = {{1'd0}, roundReg}; // @[Conditional.scala 39:67 DES_FSM.scala 53:19]
  assign pe_io_in_L = dataReg_L; // @[Conditional.scala 39:67 DES_FSM.scala 52:16]
  assign pe_io_in_R = dataReg_R; // @[Conditional.scala 39:67 DES_FSM.scala 52:16]
  assign pe_io_in_C = dataReg_C; // @[Conditional.scala 39:67 DES_FSM.scala 52:16]
  assign pe_io_in_D = dataReg_D; // @[Conditional.scala 39:67 DES_FSM.scala 52:16]
  always @(posedge clock) begin
    if (reset) begin // @[DES_FSM.scala 16:25]
      stateReg <= 3'h0; // @[DES_FSM.scala 16:25]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io_in_valid) begin // @[DES_FSM.scala 38:25]
        stateReg <= 3'h1; // @[DES_FSM.scala 41:18]
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      stateReg <= 3'h2; // @[DES_FSM.scala 49:16]
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      stateReg <= _GEN_3;
    end else begin
      stateReg <= _GEN_9;
    end
    if (reset) begin // @[DES_FSM.scala 17:25]
      roundReg <= 4'h0; // @[DES_FSM.scala 17:25]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        roundReg <= 4'h0; // @[DES_FSM.scala 48:16]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        roundReg <= _T_6; // @[DES_FSM.scala 55:16]
      end
    end
    if (reset) begin // @[DES_FSM.scala 18:24]
      textReg <= 64'h0; // @[DES_FSM.scala 18:24]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io_in_valid) begin // @[DES_FSM.scala 38:25]
        textReg <= io_in_bits_text; // @[DES_FSM.scala 39:17]
      end
    end
    if (reset) begin // @[DES_FSM.scala 19:23]
      keyReg <= 64'h0; // @[DES_FSM.scala 19:23]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io_in_valid) begin // @[DES_FSM.scala 38:25]
        keyReg <= io_in_bits_key; // @[DES_FSM.scala 40:16]
      end
    end
    if (reset) begin // @[DES_FSM.scala 20:24]
      dataReg_L <= 32'h0; // @[DES_FSM.scala 20:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_L <= ip_io_out_L; // @[DES_FSM.scala 47:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_L <= pe_io_out_L; // @[DES_FSM.scala 54:15]
      end
    end
    if (reset) begin // @[DES_FSM.scala 20:24]
      dataReg_R <= 32'h0; // @[DES_FSM.scala 20:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_R <= ip_io_out_R; // @[DES_FSM.scala 47:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_R <= pe_io_out_R; // @[DES_FSM.scala 54:15]
      end
    end
    if (reset) begin // @[DES_FSM.scala 20:24]
      dataReg_C <= 28'h0; // @[DES_FSM.scala 20:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_C <= ip_io_out_C; // @[DES_FSM.scala 47:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_C <= pe_io_out_C; // @[DES_FSM.scala 54:15]
      end
    end
    if (reset) begin // @[DES_FSM.scala 20:24]
      dataReg_D <= 28'h0; // @[DES_FSM.scala 20:24]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Conditional.scala 39:67]
        dataReg_D <= ip_io_out_D; // @[DES_FSM.scala 47:15]
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        dataReg_D <= pe_io_out_D; // @[DES_FSM.scala 54:15]
      end
    end
    if (reset) begin // @[DES_FSM.scala 21:27]
      resultsReg <= 64'h0; // @[DES_FSM.scala 21:27]
    end else if (!(_T_2)) begin // @[Conditional.scala 40:58]
      if (!(_T_3)) begin // @[Conditional.scala 39:67]
        if (!(_T_4)) begin // @[Conditional.scala 39:67]
          resultsReg <= _GEN_8;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  roundReg = _RAND_1[3:0];
  _RAND_2 = {2{`RANDOM}};
  textReg = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  keyReg = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  dataReg_L = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  dataReg_R = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  dataReg_C = _RAND_6[27:0];
  _RAND_7 = {1{`RANDOM}};
  dataReg_D = _RAND_7[27:0];
  _RAND_8 = {2{`RANDOM}};
  resultsReg = _RAND_8[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
