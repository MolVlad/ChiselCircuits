module AES_InitialOperation(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits_text,
  input  [127:0] io_in_bits_key,
  input          io_out_ready,
  output         io_out_valid,
  output [7:0]   io_out_bits_state_0_0,
  output [7:0]   io_out_bits_state_0_1,
  output [7:0]   io_out_bits_state_0_2,
  output [7:0]   io_out_bits_state_0_3,
  output [7:0]   io_out_bits_state_1_0,
  output [7:0]   io_out_bits_state_1_1,
  output [7:0]   io_out_bits_state_1_2,
  output [7:0]   io_out_bits_state_1_3,
  output [7:0]   io_out_bits_state_2_0,
  output [7:0]   io_out_bits_state_2_1,
  output [7:0]   io_out_bits_state_2_2,
  output [7:0]   io_out_bits_state_2_3,
  output [7:0]   io_out_bits_state_3_0,
  output [7:0]   io_out_bits_state_3_1,
  output [7:0]   io_out_bits_state_3_2,
  output [7:0]   io_out_bits_state_3_3,
  output [7:0]   io_out_bits_key_0_0,
  output [7:0]   io_out_bits_key_0_1,
  output [7:0]   io_out_bits_key_0_2,
  output [7:0]   io_out_bits_key_0_3,
  output [7:0]   io_out_bits_key_1_0,
  output [7:0]   io_out_bits_key_1_1,
  output [7:0]   io_out_bits_key_1_2,
  output [7:0]   io_out_bits_key_1_3,
  output [7:0]   io_out_bits_key_2_0,
  output [7:0]   io_out_bits_key_2_1,
  output [7:0]   io_out_bits_key_2_2,
  output [7:0]   io_out_bits_key_2_3,
  output [7:0]   io_out_bits_key_3_0,
  output [7:0]   io_out_bits_key_3_1,
  output [7:0]   io_out_bits_key_3_2,
  output [7:0]   io_out_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] data_0_text; // @[AES_PipelinedElasticBuffer.scala 65:21]
  reg [127:0] data_0_key; // @[AES_PipelinedElasticBuffer.scala 65:21]
  reg [127:0] data_1_text; // @[AES_PipelinedElasticBuffer.scala 65:21]
  reg [127:0] data_1_key; // @[AES_PipelinedElasticBuffer.scala 65:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 66:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 67:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 68:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 68:21]
  wire [127:0] input_text = head ? data_1_text : data_0_text; // @[AES_PipelinedElasticBuffer.scala 73:9 AES_PipelinedElasticBuffer.scala 73:9]
  wire [127:0] input_key = head ? data_1_key : data_0_key; // @[AES_PipelinedElasticBuffer.scala 73:9 AES_PipelinedElasticBuffer.scala 73:9]
  wire  _GEN_5 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 76:23 AES_PipelinedElasticBuffer.scala 76:23]
  wire  _GEN_26 = ~tail; // @[AES_PipelinedElasticBuffer.scala 77:16 AES_PipelinedElasticBuffer.scala 77:16 AES_PipelinedElasticBuffer.scala 68:21]
  wire  _GEN_6 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 77:16 AES_PipelinedElasticBuffer.scala 77:16 AES_PipelinedElasticBuffer.scala 68:21]
  wire  _GEN_7 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 77:16 AES_PipelinedElasticBuffer.scala 77:16 AES_PipelinedElasticBuffer.scala 68:21]
  wire  _GEN_12 = io_in_valid & ~_GEN_5 ? _GEN_6 : full_0; // @[AES_PipelinedElasticBuffer.scala 76:36 AES_PipelinedElasticBuffer.scala 68:21]
  wire  _GEN_13 = io_in_valid & ~_GEN_5 ? _GEN_7 : full_1; // @[AES_PipelinedElasticBuffer.scala 76:36 AES_PipelinedElasticBuffer.scala 68:21]
  wire  _GEN_20 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 83:21 AES_PipelinedElasticBuffer.scala 83:21]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 70:18]
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 71:27]
  assign io_out_bits_state_0_0 = input_text[127:120]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_0_1 = input_text[119:112]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_0_2 = input_text[111:104]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_0_3 = input_text[103:96]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_1_0 = input_text[95:88]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_1_1 = input_text[87:80]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_1_2 = input_text[79:72]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_1_3 = input_text[71:64]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_2_0 = input_text[63:56]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_2_1 = input_text[55:48]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_2_2 = input_text[47:40]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_2_3 = input_text[39:32]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_3_0 = input_text[31:24]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_3_1 = input_text[23:16]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_3_2 = input_text[15:8]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_state_3_3 = input_text[7:0]; // @[AES_PipelinedElasticBuffer.scala 91:43]
  assign io_out_bits_key_0_0 = input_key[127:120]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_0_1 = input_key[119:112]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_0_2 = input_key[111:104]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_0_3 = input_key[103:96]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_1_0 = input_key[95:88]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_1_1 = input_key[87:80]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_1_2 = input_key[79:72]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_1_3 = input_key[71:64]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_2_0 = input_key[63:56]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_2_1 = input_key[55:48]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_2_2 = input_key[47:40]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_2_3 = input_key[39:32]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_3_0 = input_key[31:24]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_3_1 = input_key[23:16]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_3_2 = input_key[15:8]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  assign io_out_bits_key_3_3 = input_key[7:0]; // @[AES_PipelinedElasticBuffer.scala 92:40]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 65:21]
      data_0_text <= 128'h0; // @[AES_PipelinedElasticBuffer.scala 65:21]
    end else if (io_in_valid & ~_GEN_5) begin // @[AES_PipelinedElasticBuffer.scala 76:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 78:16]
        data_0_text <= io_in_bits_text; // @[AES_PipelinedElasticBuffer.scala 78:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 65:21]
      data_0_key <= 128'h0; // @[AES_PipelinedElasticBuffer.scala 65:21]
    end else if (io_in_valid & ~_GEN_5) begin // @[AES_PipelinedElasticBuffer.scala 76:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 78:16]
        data_0_key <= io_in_bits_key; // @[AES_PipelinedElasticBuffer.scala 78:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 65:21]
      data_1_text <= 128'h0; // @[AES_PipelinedElasticBuffer.scala 65:21]
    end else if (io_in_valid & ~_GEN_5) begin // @[AES_PipelinedElasticBuffer.scala 76:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 78:16]
        data_1_text <= io_in_bits_text; // @[AES_PipelinedElasticBuffer.scala 78:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 65:21]
      data_1_key <= 128'h0; // @[AES_PipelinedElasticBuffer.scala 65:21]
    end else if (io_in_valid & ~_GEN_5) begin // @[AES_PipelinedElasticBuffer.scala 76:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 78:16]
        data_1_key <= io_in_bits_key; // @[AES_PipelinedElasticBuffer.scala 78:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 66:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 66:21]
    end else if (io_out_ready & _GEN_20) begin // @[AES_PipelinedElasticBuffer.scala 83:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 85:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 67:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 67:21]
    end else if (io_in_valid & ~_GEN_5) begin // @[AES_PipelinedElasticBuffer.scala 76:36]
      tail <= _GEN_26; // @[AES_PipelinedElasticBuffer.scala 79:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 68:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 68:21]
    end else if (io_out_ready & _GEN_20) begin // @[AES_PipelinedElasticBuffer.scala 83:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 84:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 84:16]
      end else begin
        full_0 <= _GEN_12;
      end
    end else begin
      full_0 <= _GEN_12;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 68:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 68:21]
    end else if (io_out_ready & _GEN_20) begin // @[AES_PipelinedElasticBuffer.scala 83:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 84:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 84:16]
      end else begin
        full_1 <= _GEN_13;
      end
    end else begin
      full_1 <= _GEN_13;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  data_0_text = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  data_0_key = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  data_1_text = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  data_1_key = _RAND_3[127:0];
  _RAND_4 = {1{`RANDOM}};
  head = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tail = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  full_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  full_1 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_FinalOperation(
  input          clock,
  input          reset,
  input          io_out_ready,
  output         io_out_valid,
  output [127:0] io_out_bits,
  output         io_in_ready,
  input          io_in_valid,
  input  [7:0]   io_in_bits_state_0_0,
  input  [7:0]   io_in_bits_state_0_1,
  input  [7:0]   io_in_bits_state_0_2,
  input  [7:0]   io_in_bits_state_0_3,
  input  [7:0]   io_in_bits_state_1_0,
  input  [7:0]   io_in_bits_state_1_1,
  input  [7:0]   io_in_bits_state_1_2,
  input  [7:0]   io_in_bits_state_1_3,
  input  [7:0]   io_in_bits_state_2_0,
  input  [7:0]   io_in_bits_state_2_1,
  input  [7:0]   io_in_bits_state_2_2,
  input  [7:0]   io_in_bits_state_2_3,
  input  [7:0]   io_in_bits_state_3_0,
  input  [7:0]   io_in_bits_state_3_1,
  input  [7:0]   io_in_bits_state_3_2,
  input  [7:0]   io_in_bits_state_3_3,
  input  [7:0]   io_in_bits_key_0_0,
  input  [7:0]   io_in_bits_key_0_1,
  input  [7:0]   io_in_bits_key_0_2,
  input  [7:0]   io_in_bits_key_0_3,
  input  [7:0]   io_in_bits_key_1_0,
  input  [7:0]   io_in_bits_key_1_1,
  input  [7:0]   io_in_bits_key_1_2,
  input  [7:0]   io_in_bits_key_1_3,
  input  [7:0]   io_in_bits_key_2_0,
  input  [7:0]   io_in_bits_key_2_1,
  input  [7:0]   io_in_bits_key_2_2,
  input  [7:0]   io_in_bits_key_2_3,
  input  [7:0]   io_in_bits_key_3_0,
  input  [7:0]   io_in_bits_key_3_1,
  input  [7:0]   io_in_bits_key_3_2,
  input  [7:0]   io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 105:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 106:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 107:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 108:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 108:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 113:9 AES_PipelinedElasticBuffer.scala 113:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 116:23 AES_PipelinedElasticBuffer.scala 116:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 117:16 AES_PipelinedElasticBuffer.scala 117:16 AES_PipelinedElasticBuffer.scala 108:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 117:16 AES_PipelinedElasticBuffer.scala 117:16 AES_PipelinedElasticBuffer.scala 108:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 117:16 AES_PipelinedElasticBuffer.scala 117:16 AES_PipelinedElasticBuffer.scala 108:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 116:36 AES_PipelinedElasticBuffer.scala 108:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 116:36 AES_PipelinedElasticBuffer.scala 108:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 123:21 AES_PipelinedElasticBuffer.scala 123:21]
  wire [7:0] hi_hi_hi_hi = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 129:34]
  wire [7:0] hi_hi_hi_lo = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 129:68]
  wire [7:0] hi_hi_lo_hi = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 130:22]
  wire [7:0] hi_hi_lo_lo = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 130:56]
  wire [7:0] hi_lo_hi_hi = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 131:22]
  wire [7:0] hi_lo_hi_lo = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 131:56]
  wire [7:0] hi_lo_lo_hi = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 132:22]
  wire [7:0] hi_lo_lo_lo = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 132:56]
  wire [7:0] lo_hi_hi_hi = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 133:22]
  wire [7:0] lo_hi_hi_lo = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 133:56]
  wire [7:0] lo_hi_lo_hi = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 134:22]
  wire [7:0] lo_hi_lo_lo = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 134:56]
  wire [7:0] lo_lo_hi_hi = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 135:22]
  wire [7:0] lo_lo_hi_lo = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 135:56]
  wire [7:0] lo_lo_lo_hi = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 136:22]
  wire [7:0] lo_lo_lo_lo = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 136:56]
  wire [63:0] lo = {lo_hi_hi_hi,lo_hi_hi_lo,lo_hi_lo_hi,lo_hi_lo_lo,lo_lo_hi_hi,lo_lo_hi_lo,lo_lo_lo_hi,lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] hi = {hi_hi_hi_hi,hi_hi_hi_lo,hi_hi_lo_hi,hi_hi_lo_lo,hi_lo_hi_hi,hi_lo_hi_lo,hi_lo_lo_hi,hi_lo_lo_lo}; // @[Cat.scala 30:58]
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 111:27]
  assign io_out_bits = {hi,lo}; // @[Cat.scala 30:58]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 110:18]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 105:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 105:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 118:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 118:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 106:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 106:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 123:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 125:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 107:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 107:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 116:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 119:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 108:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 108:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 123:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 124:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 124:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 108:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 108:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 123:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 124:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 124:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_S(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _GEN_1 = 4'h0 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h7c : 8'h63; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_2 = 4'h0 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h77 : _GEN_1; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_3 = 4'h0 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h7b : _GEN_2; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_4 = 4'h0 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hf2 : _GEN_3; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_5 = 4'h0 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h6b : _GEN_4; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_6 = 4'h0 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h6f : _GEN_5; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_7 = 4'h0 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hc5 : _GEN_6; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_8 = 4'h0 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h30 : _GEN_7; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_9 = 4'h0 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h1 : _GEN_8; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_10 = 4'h0 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h67 : _GEN_9; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_11 = 4'h0 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h2b : _GEN_10; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_12 = 4'h0 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hfe : _GEN_11; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_13 = 4'h0 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hd7 : _GEN_12; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_14 = 4'h0 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hab : _GEN_13; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_15 = 4'h0 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h76 : _GEN_14; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_16 = 4'h1 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hca : _GEN_15; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_17 = 4'h1 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h82 : _GEN_16; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_18 = 4'h1 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'hc9 : _GEN_17; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_19 = 4'h1 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h7d : _GEN_18; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_20 = 4'h1 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hfa : _GEN_19; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_21 = 4'h1 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h59 : _GEN_20; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_22 = 4'h1 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h47 : _GEN_21; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_23 = 4'h1 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hf0 : _GEN_22; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_24 = 4'h1 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'had : _GEN_23; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_25 = 4'h1 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hd4 : _GEN_24; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_26 = 4'h1 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'ha2 : _GEN_25; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_27 = 4'h1 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'haf : _GEN_26; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_28 = 4'h1 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h9c : _GEN_27; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_29 = 4'h1 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'ha4 : _GEN_28; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_30 = 4'h1 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h72 : _GEN_29; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_31 = 4'h1 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hc0 : _GEN_30; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_32 = 4'h2 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hb7 : _GEN_31; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_33 = 4'h2 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hfd : _GEN_32; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_34 = 4'h2 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h93 : _GEN_33; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_35 = 4'h2 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h26 : _GEN_34; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_36 = 4'h2 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h36 : _GEN_35; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_37 = 4'h2 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h3f : _GEN_36; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_38 = 4'h2 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hf7 : _GEN_37; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_39 = 4'h2 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hcc : _GEN_38; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_40 = 4'h2 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h34 : _GEN_39; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_41 = 4'h2 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'ha5 : _GEN_40; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_42 = 4'h2 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'he5 : _GEN_41; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_43 = 4'h2 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hf1 : _GEN_42; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_44 = 4'h2 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h71 : _GEN_43; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_45 = 4'h2 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hd8 : _GEN_44; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_46 = 4'h2 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h31 : _GEN_45; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_47 = 4'h2 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h15 : _GEN_46; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_48 = 4'h3 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h4 : _GEN_47; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_49 = 4'h3 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hc7 : _GEN_48; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_50 = 4'h3 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h23 : _GEN_49; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_51 = 4'h3 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hc3 : _GEN_50; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_52 = 4'h3 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h18 : _GEN_51; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_53 = 4'h3 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h96 : _GEN_52; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_54 = 4'h3 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h5 : _GEN_53; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_55 = 4'h3 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h9a : _GEN_54; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_56 = 4'h3 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h7 : _GEN_55; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_57 = 4'h3 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h12 : _GEN_56; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_58 = 4'h3 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h80 : _GEN_57; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_59 = 4'h3 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'he2 : _GEN_58; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_60 = 4'h3 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'heb : _GEN_59; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_61 = 4'h3 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h27 : _GEN_60; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_62 = 4'h3 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hb2 : _GEN_61; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_63 = 4'h3 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h75 : _GEN_62; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_64 = 4'h4 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h9 : _GEN_63; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_65 = 4'h4 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h83 : _GEN_64; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_66 = 4'h4 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h2c : _GEN_65; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_67 = 4'h4 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h1a : _GEN_66; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_68 = 4'h4 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h1b : _GEN_67; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_69 = 4'h4 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h6e : _GEN_68; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_70 = 4'h4 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h5a : _GEN_69; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_71 = 4'h4 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'ha0 : _GEN_70; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_72 = 4'h4 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h52 : _GEN_71; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_73 = 4'h4 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h3b : _GEN_72; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_74 = 4'h4 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hd6 : _GEN_73; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_75 = 4'h4 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hb3 : _GEN_74; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_76 = 4'h4 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h29 : _GEN_75; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_77 = 4'h4 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'he3 : _GEN_76; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_78 = 4'h4 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h2f : _GEN_77; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_79 = 4'h4 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h84 : _GEN_78; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_80 = 4'h5 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h53 : _GEN_79; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_81 = 4'h5 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hd1 : _GEN_80; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_82 = 4'h5 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h0 : _GEN_81; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_83 = 4'h5 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hed : _GEN_82; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_84 = 4'h5 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h20 : _GEN_83; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_85 = 4'h5 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hfc : _GEN_84; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_86 = 4'h5 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hb1 : _GEN_85; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_87 = 4'h5 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h5b : _GEN_86; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_88 = 4'h5 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h6a : _GEN_87; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_89 = 4'h5 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hcb : _GEN_88; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_90 = 4'h5 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hbe : _GEN_89; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_91 = 4'h5 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h39 : _GEN_90; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_92 = 4'h5 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h4a : _GEN_91; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_93 = 4'h5 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h4c : _GEN_92; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_94 = 4'h5 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h58 : _GEN_93; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_95 = 4'h5 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hcf : _GEN_94; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_96 = 4'h6 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hd0 : _GEN_95; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_97 = 4'h6 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hef : _GEN_96; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_98 = 4'h6 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'haa : _GEN_97; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_99 = 4'h6 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hfb : _GEN_98; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_100 = 4'h6 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h43 : _GEN_99; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_101 = 4'h6 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h4d : _GEN_100; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_102 = 4'h6 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h33 : _GEN_101; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_103 = 4'h6 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h85 : _GEN_102; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_104 = 4'h6 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h45 : _GEN_103; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_105 = 4'h6 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hf9 : _GEN_104; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_106 = 4'h6 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h2 : _GEN_105; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_107 = 4'h6 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h7f : _GEN_106; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_108 = 4'h6 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h50 : _GEN_107; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_109 = 4'h6 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h3c : _GEN_108; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_110 = 4'h6 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h9f : _GEN_109; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_111 = 4'h6 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'ha8 : _GEN_110; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_112 = 4'h7 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h51 : _GEN_111; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_113 = 4'h7 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'ha3 : _GEN_112; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_114 = 4'h7 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h40 : _GEN_113; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_115 = 4'h7 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h8f : _GEN_114; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_116 = 4'h7 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h92 : _GEN_115; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_117 = 4'h7 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h9d : _GEN_116; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_118 = 4'h7 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h38 : _GEN_117; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_119 = 4'h7 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hf5 : _GEN_118; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_120 = 4'h7 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hbc : _GEN_119; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_121 = 4'h7 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hb6 : _GEN_120; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_122 = 4'h7 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hda : _GEN_121; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_123 = 4'h7 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h21 : _GEN_122; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_124 = 4'h7 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h10 : _GEN_123; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_125 = 4'h7 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hff : _GEN_124; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_126 = 4'h7 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hf3 : _GEN_125; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_127 = 4'h7 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hd2 : _GEN_126; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_128 = 4'h8 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hcd : _GEN_127; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_129 = 4'h8 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hc : _GEN_128; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_130 = 4'h8 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h13 : _GEN_129; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_131 = 4'h8 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hec : _GEN_130; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_132 = 4'h8 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h5f : _GEN_131; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_133 = 4'h8 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h97 : _GEN_132; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_134 = 4'h8 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h44 : _GEN_133; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_135 = 4'h8 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h17 : _GEN_134; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_136 = 4'h8 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hc4 : _GEN_135; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_137 = 4'h8 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'ha7 : _GEN_136; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_138 = 4'h8 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h7e : _GEN_137; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_139 = 4'h8 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h3d : _GEN_138; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_140 = 4'h8 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h64 : _GEN_139; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_141 = 4'h8 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h5d : _GEN_140; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_142 = 4'h8 == io_in[7:4] & 4'he == io_in[3:0] ? 8'h19 : _GEN_141; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_143 = 4'h8 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h73 : _GEN_142; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_144 = 4'h9 == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h60 : _GEN_143; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_145 = 4'h9 == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h81 : _GEN_144; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_146 = 4'h9 == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h4f : _GEN_145; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_147 = 4'h9 == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hdc : _GEN_146; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_148 = 4'h9 == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h22 : _GEN_147; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_149 = 4'h9 == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h2a : _GEN_148; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_150 = 4'h9 == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h90 : _GEN_149; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_151 = 4'h9 == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h88 : _GEN_150; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_152 = 4'h9 == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h46 : _GEN_151; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_153 = 4'h9 == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hee : _GEN_152; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_154 = 4'h9 == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hb8 : _GEN_153; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_155 = 4'h9 == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h14 : _GEN_154; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_156 = 4'h9 == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hde : _GEN_155; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_157 = 4'h9 == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h5e : _GEN_156; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_158 = 4'h9 == io_in[7:4] & 4'he == io_in[3:0] ? 8'hb : _GEN_157; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_159 = 4'h9 == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hdb : _GEN_158; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_160 = 4'ha == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'he0 : _GEN_159; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_161 = 4'ha == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h32 : _GEN_160; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_162 = 4'ha == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h3a : _GEN_161; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_163 = 4'ha == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'ha : _GEN_162; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_164 = 4'ha == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h49 : _GEN_163; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_165 = 4'ha == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h6 : _GEN_164; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_166 = 4'ha == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h24 : _GEN_165; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_167 = 4'ha == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h5c : _GEN_166; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_168 = 4'ha == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'hc2 : _GEN_167; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_169 = 4'ha == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hd3 : _GEN_168; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_170 = 4'ha == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hac : _GEN_169; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_171 = 4'ha == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h62 : _GEN_170; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_172 = 4'ha == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h91 : _GEN_171; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_173 = 4'ha == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h95 : _GEN_172; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_174 = 4'ha == io_in[7:4] & 4'he == io_in[3:0] ? 8'he4 : _GEN_173; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_175 = 4'ha == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h79 : _GEN_174; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_176 = 4'hb == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'he7 : _GEN_175; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_177 = 4'hb == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hc8 : _GEN_176; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_178 = 4'hb == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h37 : _GEN_177; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_179 = 4'hb == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h6d : _GEN_178; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_180 = 4'hb == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h8d : _GEN_179; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_181 = 4'hb == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hd5 : _GEN_180; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_182 = 4'hb == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h4e : _GEN_181; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_183 = 4'hb == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'ha9 : _GEN_182; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_184 = 4'hb == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h6c : _GEN_183; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_185 = 4'hb == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h56 : _GEN_184; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_186 = 4'hb == io_in[7:4] & 4'ha == io_in[3:0] ? 8'hf4 : _GEN_185; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_187 = 4'hb == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hea : _GEN_186; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_188 = 4'hb == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h65 : _GEN_187; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_189 = 4'hb == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h7a : _GEN_188; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_190 = 4'hb == io_in[7:4] & 4'he == io_in[3:0] ? 8'hae : _GEN_189; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_191 = 4'hb == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h8 : _GEN_190; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_192 = 4'hc == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'hba : _GEN_191; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_193 = 4'hc == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h78 : _GEN_192; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_194 = 4'hc == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h25 : _GEN_193; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_195 = 4'hc == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h2e : _GEN_194; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_196 = 4'hc == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h1c : _GEN_195; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_197 = 4'hc == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'ha6 : _GEN_196; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_198 = 4'hc == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hb4 : _GEN_197; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_199 = 4'hc == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'hc6 : _GEN_198; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_200 = 4'hc == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'he8 : _GEN_199; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_201 = 4'hc == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'hdd : _GEN_200; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_202 = 4'hc == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h74 : _GEN_201; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_203 = 4'hc == io_in[7:4] & 4'hb == io_in[3:0] ? 8'h1f : _GEN_202; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_204 = 4'hc == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h4b : _GEN_203; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_205 = 4'hc == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hbd : _GEN_204; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_206 = 4'hc == io_in[7:4] & 4'he == io_in[3:0] ? 8'h8b : _GEN_205; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_207 = 4'hc == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h8a : _GEN_206; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_208 = 4'hd == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h70 : _GEN_207; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_209 = 4'hd == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'h3e : _GEN_208; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_210 = 4'hd == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'hb5 : _GEN_209; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_211 = 4'hd == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h66 : _GEN_210; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_212 = 4'hd == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h48 : _GEN_211; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_213 = 4'hd == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'h3 : _GEN_212; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_214 = 4'hd == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'hf6 : _GEN_213; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_215 = 4'hd == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'he : _GEN_214; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_216 = 4'hd == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h61 : _GEN_215; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_217 = 4'hd == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h35 : _GEN_216; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_218 = 4'hd == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h57 : _GEN_217; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_219 = 4'hd == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hb9 : _GEN_218; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_220 = 4'hd == io_in[7:4] & 4'hc == io_in[3:0] ? 8'h86 : _GEN_219; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_221 = 4'hd == io_in[7:4] & 4'hd == io_in[3:0] ? 8'hc1 : _GEN_220; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_222 = 4'hd == io_in[7:4] & 4'he == io_in[3:0] ? 8'h1d : _GEN_221; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_223 = 4'hd == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h9e : _GEN_222; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_224 = 4'he == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'he1 : _GEN_223; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_225 = 4'he == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'hf8 : _GEN_224; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_226 = 4'he == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h98 : _GEN_225; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_227 = 4'he == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'h11 : _GEN_226; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_228 = 4'he == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'h69 : _GEN_227; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_229 = 4'he == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'hd9 : _GEN_228; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_230 = 4'he == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h8e : _GEN_229; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_231 = 4'he == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h94 : _GEN_230; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_232 = 4'he == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h9b : _GEN_231; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_233 = 4'he == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h1e : _GEN_232; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_234 = 4'he == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h87 : _GEN_233; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_235 = 4'he == io_in[7:4] & 4'hb == io_in[3:0] ? 8'he9 : _GEN_234; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_236 = 4'he == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hce : _GEN_235; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_237 = 4'he == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h55 : _GEN_236; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_238 = 4'he == io_in[7:4] & 4'he == io_in[3:0] ? 8'h28 : _GEN_237; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_239 = 4'he == io_in[7:4] & 4'hf == io_in[3:0] ? 8'hdf : _GEN_238; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_240 = 4'hf == io_in[7:4] & 4'h0 == io_in[3:0] ? 8'h8c : _GEN_239; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_241 = 4'hf == io_in[7:4] & 4'h1 == io_in[3:0] ? 8'ha1 : _GEN_240; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_242 = 4'hf == io_in[7:4] & 4'h2 == io_in[3:0] ? 8'h89 : _GEN_241; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_243 = 4'hf == io_in[7:4] & 4'h3 == io_in[3:0] ? 8'hd : _GEN_242; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_244 = 4'hf == io_in[7:4] & 4'h4 == io_in[3:0] ? 8'hbf : _GEN_243; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_245 = 4'hf == io_in[7:4] & 4'h5 == io_in[3:0] ? 8'he6 : _GEN_244; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_246 = 4'hf == io_in[7:4] & 4'h6 == io_in[3:0] ? 8'h42 : _GEN_245; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_247 = 4'hf == io_in[7:4] & 4'h7 == io_in[3:0] ? 8'h68 : _GEN_246; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_248 = 4'hf == io_in[7:4] & 4'h8 == io_in[3:0] ? 8'h41 : _GEN_247; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_249 = 4'hf == io_in[7:4] & 4'h9 == io_in[3:0] ? 8'h99 : _GEN_248; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_250 = 4'hf == io_in[7:4] & 4'ha == io_in[3:0] ? 8'h2d : _GEN_249; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_251 = 4'hf == io_in[7:4] & 4'hb == io_in[3:0] ? 8'hf : _GEN_250; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_252 = 4'hf == io_in[7:4] & 4'hc == io_in[3:0] ? 8'hb0 : _GEN_251; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_253 = 4'hf == io_in[7:4] & 4'hd == io_in[3:0] ? 8'h54 : _GEN_252; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  wire [7:0] _GEN_254 = 4'hf == io_in[7:4] & 4'he == io_in[3:0] ? 8'hbb : _GEN_253; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
  assign io_out = 4'hf == io_in[7:4] & 4'hf == io_in[3:0] ? 8'h16 : _GEN_254; // @[AES_PipelinedElasticBuffer.scala 426:10 AES_PipelinedElasticBuffer.scala 426:10]
endmodule
module AES_SubBytes(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3
);
  wire [7:0] PEs_0_0_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_0_0_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_0_1_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_0_1_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_0_2_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_0_2_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_0_3_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_0_3_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_1_0_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_1_0_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_1_1_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_1_1_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_1_2_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_1_2_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_1_3_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_1_3_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_2_0_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_2_0_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_2_1_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_2_1_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_2_2_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_2_2_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_2_3_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_2_3_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_3_0_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_3_0_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_3_1_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_3_1_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_3_2_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_3_2_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_3_3_io_in; // @[AES_PipelinedElasticBuffer.scala 373:22]
  wire [7:0] PEs_3_3_io_out; // @[AES_PipelinedElasticBuffer.scala 373:22]
  AES_S PEs_0_0 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_0_0_io_in),
    .io_out(PEs_0_0_io_out)
  );
  AES_S PEs_0_1 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_0_1_io_in),
    .io_out(PEs_0_1_io_out)
  );
  AES_S PEs_0_2 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_0_2_io_in),
    .io_out(PEs_0_2_io_out)
  );
  AES_S PEs_0_3 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_0_3_io_in),
    .io_out(PEs_0_3_io_out)
  );
  AES_S PEs_1_0 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_1_0_io_in),
    .io_out(PEs_1_0_io_out)
  );
  AES_S PEs_1_1 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_1_1_io_in),
    .io_out(PEs_1_1_io_out)
  );
  AES_S PEs_1_2 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_1_2_io_in),
    .io_out(PEs_1_2_io_out)
  );
  AES_S PEs_1_3 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_1_3_io_in),
    .io_out(PEs_1_3_io_out)
  );
  AES_S PEs_2_0 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_2_0_io_in),
    .io_out(PEs_2_0_io_out)
  );
  AES_S PEs_2_1 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_2_1_io_in),
    .io_out(PEs_2_1_io_out)
  );
  AES_S PEs_2_2 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_2_2_io_in),
    .io_out(PEs_2_2_io_out)
  );
  AES_S PEs_2_3 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_2_3_io_in),
    .io_out(PEs_2_3_io_out)
  );
  AES_S PEs_3_0 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_3_0_io_in),
    .io_out(PEs_3_0_io_out)
  );
  AES_S PEs_3_1 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_3_1_io_in),
    .io_out(PEs_3_1_io_out)
  );
  AES_S PEs_3_2 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_3_2_io_in),
    .io_out(PEs_3_2_io_out)
  );
  AES_S PEs_3_3 ( // @[AES_PipelinedElasticBuffer.scala 373:22]
    .io_in(PEs_3_3_io_in),
    .io_out(PEs_3_3_io_out)
  );
  assign io_out_state_0_0 = PEs_0_0_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_0_1 = PEs_0_1_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_0_2 = PEs_0_2_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_0_3 = PEs_0_3_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_1_0 = PEs_1_0_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_1_1 = PEs_1_1_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_1_2 = PEs_1_2_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_1_3 = PEs_1_3_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_2_0 = PEs_2_0_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_2_1 = PEs_2_1_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_2_2 = PEs_2_2_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_2_3 = PEs_2_3_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_3_0 = PEs_3_0_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_3_1 = PEs_3_1_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_3_2 = PEs_3_2_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign io_out_state_3_3 = PEs_3_3_io_out; // @[AES_PipelinedElasticBuffer.scala 382:26]
  assign PEs_0_0_io_in = io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_0_1_io_in = io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_0_2_io_in = io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_0_3_io_in = io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_1_0_io_in = io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_1_1_io_in = io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_1_2_io_in = io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_1_3_io_in = io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_2_0_io_in = io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_2_1_io_in = io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_2_2_io_in = io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_2_3_io_in = io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_3_0_io_in = io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_3_1_io_in = io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_3_2_io_in = io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 381:23]
  assign PEs_3_3_io_in = io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 381:23]
endmodule
module AES_ShiftRows(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3
);
  assign io_out_state_0_0 = io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 342:22]
  assign io_out_state_0_1 = io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 347:22]
  assign io_out_state_0_2 = io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 352:22]
  assign io_out_state_0_3 = io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 357:22]
  assign io_out_state_1_0 = io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 343:22]
  assign io_out_state_1_1 = io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 348:22]
  assign io_out_state_1_2 = io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 353:22]
  assign io_out_state_1_3 = io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 358:22]
  assign io_out_state_2_0 = io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 344:22]
  assign io_out_state_2_1 = io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 349:22]
  assign io_out_state_2_2 = io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 354:22]
  assign io_out_state_2_3 = io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 359:22]
  assign io_out_state_3_0 = io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 345:22]
  assign io_out_state_3_1 = io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 350:22]
  assign io_out_state_3_2 = io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 355:22]
  assign io_out_state_3_3 = io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 360:22]
endmodule
module AES_MixColumn(
  input  [7:0] io_in_0,
  input  [7:0] io_in_1,
  input  [7:0] io_in_2,
  input  [7:0] io_in_3,
  output [7:0] io_out_0,
  output [7:0] io_out_1,
  output [7:0] io_out_2,
  output [7:0] io_out_3
);
  wire [7:0] _GEN_1 = 8'h1 == io_in_0 ? 8'h2 : 8'h0; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_2 = 8'h2 == io_in_0 ? 8'h4 : _GEN_1; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_3 = 8'h3 == io_in_0 ? 8'h6 : _GEN_2; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_4 = 8'h4 == io_in_0 ? 8'h8 : _GEN_3; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_5 = 8'h5 == io_in_0 ? 8'ha : _GEN_4; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_6 = 8'h6 == io_in_0 ? 8'hc : _GEN_5; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_7 = 8'h7 == io_in_0 ? 8'he : _GEN_6; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_8 = 8'h8 == io_in_0 ? 8'h10 : _GEN_7; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_9 = 8'h9 == io_in_0 ? 8'h12 : _GEN_8; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_10 = 8'ha == io_in_0 ? 8'h14 : _GEN_9; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_11 = 8'hb == io_in_0 ? 8'h16 : _GEN_10; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_12 = 8'hc == io_in_0 ? 8'h18 : _GEN_11; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_13 = 8'hd == io_in_0 ? 8'h1a : _GEN_12; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_14 = 8'he == io_in_0 ? 8'h1c : _GEN_13; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_15 = 8'hf == io_in_0 ? 8'h1e : _GEN_14; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_16 = 8'h10 == io_in_0 ? 8'h20 : _GEN_15; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_17 = 8'h11 == io_in_0 ? 8'h22 : _GEN_16; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_18 = 8'h12 == io_in_0 ? 8'h24 : _GEN_17; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_19 = 8'h13 == io_in_0 ? 8'h26 : _GEN_18; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_20 = 8'h14 == io_in_0 ? 8'h28 : _GEN_19; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_21 = 8'h15 == io_in_0 ? 8'h2a : _GEN_20; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_22 = 8'h16 == io_in_0 ? 8'h2c : _GEN_21; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_23 = 8'h17 == io_in_0 ? 8'h2e : _GEN_22; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_24 = 8'h18 == io_in_0 ? 8'h30 : _GEN_23; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_25 = 8'h19 == io_in_0 ? 8'h32 : _GEN_24; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_26 = 8'h1a == io_in_0 ? 8'h34 : _GEN_25; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_27 = 8'h1b == io_in_0 ? 8'h36 : _GEN_26; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_28 = 8'h1c == io_in_0 ? 8'h38 : _GEN_27; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_29 = 8'h1d == io_in_0 ? 8'h3a : _GEN_28; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_30 = 8'h1e == io_in_0 ? 8'h3c : _GEN_29; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_31 = 8'h1f == io_in_0 ? 8'h3e : _GEN_30; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_32 = 8'h20 == io_in_0 ? 8'h40 : _GEN_31; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_33 = 8'h21 == io_in_0 ? 8'h42 : _GEN_32; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_34 = 8'h22 == io_in_0 ? 8'h44 : _GEN_33; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_35 = 8'h23 == io_in_0 ? 8'h46 : _GEN_34; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_36 = 8'h24 == io_in_0 ? 8'h48 : _GEN_35; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_37 = 8'h25 == io_in_0 ? 8'h4a : _GEN_36; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_38 = 8'h26 == io_in_0 ? 8'h4c : _GEN_37; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_39 = 8'h27 == io_in_0 ? 8'h4e : _GEN_38; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_40 = 8'h28 == io_in_0 ? 8'h50 : _GEN_39; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_41 = 8'h29 == io_in_0 ? 8'h52 : _GEN_40; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_42 = 8'h2a == io_in_0 ? 8'h54 : _GEN_41; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_43 = 8'h2b == io_in_0 ? 8'h56 : _GEN_42; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_44 = 8'h2c == io_in_0 ? 8'h58 : _GEN_43; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_45 = 8'h2d == io_in_0 ? 8'h5a : _GEN_44; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_46 = 8'h2e == io_in_0 ? 8'h5c : _GEN_45; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_47 = 8'h2f == io_in_0 ? 8'h5e : _GEN_46; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_48 = 8'h30 == io_in_0 ? 8'h60 : _GEN_47; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_49 = 8'h31 == io_in_0 ? 8'h62 : _GEN_48; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_50 = 8'h32 == io_in_0 ? 8'h64 : _GEN_49; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_51 = 8'h33 == io_in_0 ? 8'h66 : _GEN_50; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_52 = 8'h34 == io_in_0 ? 8'h68 : _GEN_51; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_53 = 8'h35 == io_in_0 ? 8'h6a : _GEN_52; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_54 = 8'h36 == io_in_0 ? 8'h6c : _GEN_53; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_55 = 8'h37 == io_in_0 ? 8'h6e : _GEN_54; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_56 = 8'h38 == io_in_0 ? 8'h70 : _GEN_55; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_57 = 8'h39 == io_in_0 ? 8'h72 : _GEN_56; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_58 = 8'h3a == io_in_0 ? 8'h74 : _GEN_57; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_59 = 8'h3b == io_in_0 ? 8'h76 : _GEN_58; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_60 = 8'h3c == io_in_0 ? 8'h78 : _GEN_59; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_61 = 8'h3d == io_in_0 ? 8'h7a : _GEN_60; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_62 = 8'h3e == io_in_0 ? 8'h7c : _GEN_61; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_63 = 8'h3f == io_in_0 ? 8'h7e : _GEN_62; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_64 = 8'h40 == io_in_0 ? 8'h80 : _GEN_63; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_65 = 8'h41 == io_in_0 ? 8'h82 : _GEN_64; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_66 = 8'h42 == io_in_0 ? 8'h84 : _GEN_65; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_67 = 8'h43 == io_in_0 ? 8'h86 : _GEN_66; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_68 = 8'h44 == io_in_0 ? 8'h88 : _GEN_67; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_69 = 8'h45 == io_in_0 ? 8'h8a : _GEN_68; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_70 = 8'h46 == io_in_0 ? 8'h8c : _GEN_69; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_71 = 8'h47 == io_in_0 ? 8'h8e : _GEN_70; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_72 = 8'h48 == io_in_0 ? 8'h90 : _GEN_71; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_73 = 8'h49 == io_in_0 ? 8'h92 : _GEN_72; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_74 = 8'h4a == io_in_0 ? 8'h94 : _GEN_73; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_75 = 8'h4b == io_in_0 ? 8'h96 : _GEN_74; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_76 = 8'h4c == io_in_0 ? 8'h98 : _GEN_75; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_77 = 8'h4d == io_in_0 ? 8'h9a : _GEN_76; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_78 = 8'h4e == io_in_0 ? 8'h9c : _GEN_77; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_79 = 8'h4f == io_in_0 ? 8'h9e : _GEN_78; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_80 = 8'h50 == io_in_0 ? 8'ha0 : _GEN_79; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_81 = 8'h51 == io_in_0 ? 8'ha2 : _GEN_80; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_82 = 8'h52 == io_in_0 ? 8'ha4 : _GEN_81; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_83 = 8'h53 == io_in_0 ? 8'ha6 : _GEN_82; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_84 = 8'h54 == io_in_0 ? 8'ha8 : _GEN_83; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_85 = 8'h55 == io_in_0 ? 8'haa : _GEN_84; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_86 = 8'h56 == io_in_0 ? 8'hac : _GEN_85; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_87 = 8'h57 == io_in_0 ? 8'hae : _GEN_86; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_88 = 8'h58 == io_in_0 ? 8'hb0 : _GEN_87; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_89 = 8'h59 == io_in_0 ? 8'hb2 : _GEN_88; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_90 = 8'h5a == io_in_0 ? 8'hb4 : _GEN_89; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_91 = 8'h5b == io_in_0 ? 8'hb6 : _GEN_90; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_92 = 8'h5c == io_in_0 ? 8'hb8 : _GEN_91; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_93 = 8'h5d == io_in_0 ? 8'hba : _GEN_92; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_94 = 8'h5e == io_in_0 ? 8'hbc : _GEN_93; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_95 = 8'h5f == io_in_0 ? 8'hbe : _GEN_94; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_96 = 8'h60 == io_in_0 ? 8'hc0 : _GEN_95; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_97 = 8'h61 == io_in_0 ? 8'hc2 : _GEN_96; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_98 = 8'h62 == io_in_0 ? 8'hc4 : _GEN_97; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_99 = 8'h63 == io_in_0 ? 8'hc6 : _GEN_98; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_100 = 8'h64 == io_in_0 ? 8'hc8 : _GEN_99; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_101 = 8'h65 == io_in_0 ? 8'hca : _GEN_100; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_102 = 8'h66 == io_in_0 ? 8'hcc : _GEN_101; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_103 = 8'h67 == io_in_0 ? 8'hce : _GEN_102; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_104 = 8'h68 == io_in_0 ? 8'hd0 : _GEN_103; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_105 = 8'h69 == io_in_0 ? 8'hd2 : _GEN_104; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_106 = 8'h6a == io_in_0 ? 8'hd4 : _GEN_105; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_107 = 8'h6b == io_in_0 ? 8'hd6 : _GEN_106; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_108 = 8'h6c == io_in_0 ? 8'hd8 : _GEN_107; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_109 = 8'h6d == io_in_0 ? 8'hda : _GEN_108; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_110 = 8'h6e == io_in_0 ? 8'hdc : _GEN_109; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_111 = 8'h6f == io_in_0 ? 8'hde : _GEN_110; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_112 = 8'h70 == io_in_0 ? 8'he0 : _GEN_111; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_113 = 8'h71 == io_in_0 ? 8'he2 : _GEN_112; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_114 = 8'h72 == io_in_0 ? 8'he4 : _GEN_113; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_115 = 8'h73 == io_in_0 ? 8'he6 : _GEN_114; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_116 = 8'h74 == io_in_0 ? 8'he8 : _GEN_115; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_117 = 8'h75 == io_in_0 ? 8'hea : _GEN_116; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_118 = 8'h76 == io_in_0 ? 8'hec : _GEN_117; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_119 = 8'h77 == io_in_0 ? 8'hee : _GEN_118; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_120 = 8'h78 == io_in_0 ? 8'hf0 : _GEN_119; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_121 = 8'h79 == io_in_0 ? 8'hf2 : _GEN_120; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_122 = 8'h7a == io_in_0 ? 8'hf4 : _GEN_121; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_123 = 8'h7b == io_in_0 ? 8'hf6 : _GEN_122; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_124 = 8'h7c == io_in_0 ? 8'hf8 : _GEN_123; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_125 = 8'h7d == io_in_0 ? 8'hfa : _GEN_124; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_126 = 8'h7e == io_in_0 ? 8'hfc : _GEN_125; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_127 = 8'h7f == io_in_0 ? 8'hfe : _GEN_126; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_128 = 8'h80 == io_in_0 ? 8'h1b : _GEN_127; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_129 = 8'h81 == io_in_0 ? 8'h19 : _GEN_128; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_130 = 8'h82 == io_in_0 ? 8'h1f : _GEN_129; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_131 = 8'h83 == io_in_0 ? 8'h1d : _GEN_130; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_132 = 8'h84 == io_in_0 ? 8'h13 : _GEN_131; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_133 = 8'h85 == io_in_0 ? 8'h11 : _GEN_132; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_134 = 8'h86 == io_in_0 ? 8'h17 : _GEN_133; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_135 = 8'h87 == io_in_0 ? 8'h15 : _GEN_134; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_136 = 8'h88 == io_in_0 ? 8'hb : _GEN_135; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_137 = 8'h89 == io_in_0 ? 8'h9 : _GEN_136; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_138 = 8'h8a == io_in_0 ? 8'hf : _GEN_137; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_139 = 8'h8b == io_in_0 ? 8'hd : _GEN_138; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_140 = 8'h8c == io_in_0 ? 8'h3 : _GEN_139; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_141 = 8'h8d == io_in_0 ? 8'h1 : _GEN_140; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_142 = 8'h8e == io_in_0 ? 8'h7 : _GEN_141; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_143 = 8'h8f == io_in_0 ? 8'h5 : _GEN_142; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_144 = 8'h90 == io_in_0 ? 8'h3b : _GEN_143; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_145 = 8'h91 == io_in_0 ? 8'h39 : _GEN_144; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_146 = 8'h92 == io_in_0 ? 8'h3f : _GEN_145; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_147 = 8'h93 == io_in_0 ? 8'h3d : _GEN_146; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_148 = 8'h94 == io_in_0 ? 8'h33 : _GEN_147; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_149 = 8'h95 == io_in_0 ? 8'h31 : _GEN_148; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_150 = 8'h96 == io_in_0 ? 8'h37 : _GEN_149; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_151 = 8'h97 == io_in_0 ? 8'h35 : _GEN_150; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_152 = 8'h98 == io_in_0 ? 8'h2b : _GEN_151; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_153 = 8'h99 == io_in_0 ? 8'h29 : _GEN_152; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_154 = 8'h9a == io_in_0 ? 8'h2f : _GEN_153; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_155 = 8'h9b == io_in_0 ? 8'h2d : _GEN_154; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_156 = 8'h9c == io_in_0 ? 8'h23 : _GEN_155; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_157 = 8'h9d == io_in_0 ? 8'h21 : _GEN_156; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_158 = 8'h9e == io_in_0 ? 8'h27 : _GEN_157; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_159 = 8'h9f == io_in_0 ? 8'h25 : _GEN_158; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_160 = 8'ha0 == io_in_0 ? 8'h5b : _GEN_159; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_161 = 8'ha1 == io_in_0 ? 8'h59 : _GEN_160; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_162 = 8'ha2 == io_in_0 ? 8'h5f : _GEN_161; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_163 = 8'ha3 == io_in_0 ? 8'h5d : _GEN_162; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_164 = 8'ha4 == io_in_0 ? 8'h53 : _GEN_163; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_165 = 8'ha5 == io_in_0 ? 8'h51 : _GEN_164; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_166 = 8'ha6 == io_in_0 ? 8'h57 : _GEN_165; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_167 = 8'ha7 == io_in_0 ? 8'h55 : _GEN_166; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_168 = 8'ha8 == io_in_0 ? 8'h4b : _GEN_167; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_169 = 8'ha9 == io_in_0 ? 8'h49 : _GEN_168; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_170 = 8'haa == io_in_0 ? 8'h4f : _GEN_169; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_171 = 8'hab == io_in_0 ? 8'h4d : _GEN_170; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_172 = 8'hac == io_in_0 ? 8'h43 : _GEN_171; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_173 = 8'had == io_in_0 ? 8'h41 : _GEN_172; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_174 = 8'hae == io_in_0 ? 8'h47 : _GEN_173; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_175 = 8'haf == io_in_0 ? 8'h45 : _GEN_174; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_176 = 8'hb0 == io_in_0 ? 8'h7b : _GEN_175; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_177 = 8'hb1 == io_in_0 ? 8'h79 : _GEN_176; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_178 = 8'hb2 == io_in_0 ? 8'h7f : _GEN_177; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_179 = 8'hb3 == io_in_0 ? 8'h7d : _GEN_178; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_180 = 8'hb4 == io_in_0 ? 8'h73 : _GEN_179; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_181 = 8'hb5 == io_in_0 ? 8'h71 : _GEN_180; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_182 = 8'hb6 == io_in_0 ? 8'h77 : _GEN_181; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_183 = 8'hb7 == io_in_0 ? 8'h75 : _GEN_182; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_184 = 8'hb8 == io_in_0 ? 8'h6b : _GEN_183; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_185 = 8'hb9 == io_in_0 ? 8'h69 : _GEN_184; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_186 = 8'hba == io_in_0 ? 8'h6f : _GEN_185; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_187 = 8'hbb == io_in_0 ? 8'h6d : _GEN_186; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_188 = 8'hbc == io_in_0 ? 8'h63 : _GEN_187; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_189 = 8'hbd == io_in_0 ? 8'h61 : _GEN_188; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_190 = 8'hbe == io_in_0 ? 8'h67 : _GEN_189; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_191 = 8'hbf == io_in_0 ? 8'h65 : _GEN_190; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_192 = 8'hc0 == io_in_0 ? 8'h9b : _GEN_191; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_193 = 8'hc1 == io_in_0 ? 8'h99 : _GEN_192; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_194 = 8'hc2 == io_in_0 ? 8'h9f : _GEN_193; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_195 = 8'hc3 == io_in_0 ? 8'h9d : _GEN_194; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_196 = 8'hc4 == io_in_0 ? 8'h93 : _GEN_195; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_197 = 8'hc5 == io_in_0 ? 8'h91 : _GEN_196; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_198 = 8'hc6 == io_in_0 ? 8'h97 : _GEN_197; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_199 = 8'hc7 == io_in_0 ? 8'h95 : _GEN_198; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_200 = 8'hc8 == io_in_0 ? 8'h8b : _GEN_199; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_201 = 8'hc9 == io_in_0 ? 8'h89 : _GEN_200; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_202 = 8'hca == io_in_0 ? 8'h8f : _GEN_201; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_203 = 8'hcb == io_in_0 ? 8'h8d : _GEN_202; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_204 = 8'hcc == io_in_0 ? 8'h83 : _GEN_203; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_205 = 8'hcd == io_in_0 ? 8'h81 : _GEN_204; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_206 = 8'hce == io_in_0 ? 8'h87 : _GEN_205; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_207 = 8'hcf == io_in_0 ? 8'h85 : _GEN_206; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_208 = 8'hd0 == io_in_0 ? 8'hbb : _GEN_207; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_209 = 8'hd1 == io_in_0 ? 8'hb9 : _GEN_208; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_210 = 8'hd2 == io_in_0 ? 8'hbf : _GEN_209; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_211 = 8'hd3 == io_in_0 ? 8'hbd : _GEN_210; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_212 = 8'hd4 == io_in_0 ? 8'hb3 : _GEN_211; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_213 = 8'hd5 == io_in_0 ? 8'hb1 : _GEN_212; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_214 = 8'hd6 == io_in_0 ? 8'hb7 : _GEN_213; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_215 = 8'hd7 == io_in_0 ? 8'hb5 : _GEN_214; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_216 = 8'hd8 == io_in_0 ? 8'hab : _GEN_215; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_217 = 8'hd9 == io_in_0 ? 8'ha9 : _GEN_216; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_218 = 8'hda == io_in_0 ? 8'haf : _GEN_217; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_219 = 8'hdb == io_in_0 ? 8'had : _GEN_218; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_220 = 8'hdc == io_in_0 ? 8'ha3 : _GEN_219; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_221 = 8'hdd == io_in_0 ? 8'ha1 : _GEN_220; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_222 = 8'hde == io_in_0 ? 8'ha7 : _GEN_221; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_223 = 8'hdf == io_in_0 ? 8'ha5 : _GEN_222; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_224 = 8'he0 == io_in_0 ? 8'hdb : _GEN_223; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_225 = 8'he1 == io_in_0 ? 8'hd9 : _GEN_224; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_226 = 8'he2 == io_in_0 ? 8'hdf : _GEN_225; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_227 = 8'he3 == io_in_0 ? 8'hdd : _GEN_226; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_228 = 8'he4 == io_in_0 ? 8'hd3 : _GEN_227; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_229 = 8'he5 == io_in_0 ? 8'hd1 : _GEN_228; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_230 = 8'he6 == io_in_0 ? 8'hd7 : _GEN_229; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_231 = 8'he7 == io_in_0 ? 8'hd5 : _GEN_230; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_232 = 8'he8 == io_in_0 ? 8'hcb : _GEN_231; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_233 = 8'he9 == io_in_0 ? 8'hc9 : _GEN_232; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_234 = 8'hea == io_in_0 ? 8'hcf : _GEN_233; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_235 = 8'heb == io_in_0 ? 8'hcd : _GEN_234; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_236 = 8'hec == io_in_0 ? 8'hc3 : _GEN_235; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_237 = 8'hed == io_in_0 ? 8'hc1 : _GEN_236; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_238 = 8'hee == io_in_0 ? 8'hc7 : _GEN_237; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_239 = 8'hef == io_in_0 ? 8'hc5 : _GEN_238; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_240 = 8'hf0 == io_in_0 ? 8'hfb : _GEN_239; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_241 = 8'hf1 == io_in_0 ? 8'hf9 : _GEN_240; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_242 = 8'hf2 == io_in_0 ? 8'hff : _GEN_241; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_243 = 8'hf3 == io_in_0 ? 8'hfd : _GEN_242; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_244 = 8'hf4 == io_in_0 ? 8'hf3 : _GEN_243; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_245 = 8'hf5 == io_in_0 ? 8'hf1 : _GEN_244; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_246 = 8'hf6 == io_in_0 ? 8'hf7 : _GEN_245; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_247 = 8'hf7 == io_in_0 ? 8'hf5 : _GEN_246; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_248 = 8'hf8 == io_in_0 ? 8'heb : _GEN_247; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_249 = 8'hf9 == io_in_0 ? 8'he9 : _GEN_248; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_250 = 8'hfa == io_in_0 ? 8'hef : _GEN_249; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_251 = 8'hfb == io_in_0 ? 8'hed : _GEN_250; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_252 = 8'hfc == io_in_0 ? 8'he3 : _GEN_251; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_253 = 8'hfd == io_in_0 ? 8'he1 : _GEN_252; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_254 = 8'hfe == io_in_0 ? 8'he7 : _GEN_253; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_255 = 8'hff == io_in_0 ? 8'he5 : _GEN_254; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_257 = 8'h1 == io_in_1 ? 8'h2 : 8'h0; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_258 = 8'h2 == io_in_1 ? 8'h4 : _GEN_257; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_259 = 8'h3 == io_in_1 ? 8'h6 : _GEN_258; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_260 = 8'h4 == io_in_1 ? 8'h8 : _GEN_259; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_261 = 8'h5 == io_in_1 ? 8'ha : _GEN_260; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_262 = 8'h6 == io_in_1 ? 8'hc : _GEN_261; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_263 = 8'h7 == io_in_1 ? 8'he : _GEN_262; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_264 = 8'h8 == io_in_1 ? 8'h10 : _GEN_263; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_265 = 8'h9 == io_in_1 ? 8'h12 : _GEN_264; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_266 = 8'ha == io_in_1 ? 8'h14 : _GEN_265; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_267 = 8'hb == io_in_1 ? 8'h16 : _GEN_266; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_268 = 8'hc == io_in_1 ? 8'h18 : _GEN_267; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_269 = 8'hd == io_in_1 ? 8'h1a : _GEN_268; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_270 = 8'he == io_in_1 ? 8'h1c : _GEN_269; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_271 = 8'hf == io_in_1 ? 8'h1e : _GEN_270; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_272 = 8'h10 == io_in_1 ? 8'h20 : _GEN_271; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_273 = 8'h11 == io_in_1 ? 8'h22 : _GEN_272; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_274 = 8'h12 == io_in_1 ? 8'h24 : _GEN_273; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_275 = 8'h13 == io_in_1 ? 8'h26 : _GEN_274; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_276 = 8'h14 == io_in_1 ? 8'h28 : _GEN_275; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_277 = 8'h15 == io_in_1 ? 8'h2a : _GEN_276; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_278 = 8'h16 == io_in_1 ? 8'h2c : _GEN_277; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_279 = 8'h17 == io_in_1 ? 8'h2e : _GEN_278; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_280 = 8'h18 == io_in_1 ? 8'h30 : _GEN_279; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_281 = 8'h19 == io_in_1 ? 8'h32 : _GEN_280; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_282 = 8'h1a == io_in_1 ? 8'h34 : _GEN_281; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_283 = 8'h1b == io_in_1 ? 8'h36 : _GEN_282; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_284 = 8'h1c == io_in_1 ? 8'h38 : _GEN_283; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_285 = 8'h1d == io_in_1 ? 8'h3a : _GEN_284; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_286 = 8'h1e == io_in_1 ? 8'h3c : _GEN_285; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_287 = 8'h1f == io_in_1 ? 8'h3e : _GEN_286; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_288 = 8'h20 == io_in_1 ? 8'h40 : _GEN_287; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_289 = 8'h21 == io_in_1 ? 8'h42 : _GEN_288; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_290 = 8'h22 == io_in_1 ? 8'h44 : _GEN_289; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_291 = 8'h23 == io_in_1 ? 8'h46 : _GEN_290; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_292 = 8'h24 == io_in_1 ? 8'h48 : _GEN_291; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_293 = 8'h25 == io_in_1 ? 8'h4a : _GEN_292; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_294 = 8'h26 == io_in_1 ? 8'h4c : _GEN_293; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_295 = 8'h27 == io_in_1 ? 8'h4e : _GEN_294; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_296 = 8'h28 == io_in_1 ? 8'h50 : _GEN_295; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_297 = 8'h29 == io_in_1 ? 8'h52 : _GEN_296; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_298 = 8'h2a == io_in_1 ? 8'h54 : _GEN_297; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_299 = 8'h2b == io_in_1 ? 8'h56 : _GEN_298; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_300 = 8'h2c == io_in_1 ? 8'h58 : _GEN_299; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_301 = 8'h2d == io_in_1 ? 8'h5a : _GEN_300; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_302 = 8'h2e == io_in_1 ? 8'h5c : _GEN_301; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_303 = 8'h2f == io_in_1 ? 8'h5e : _GEN_302; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_304 = 8'h30 == io_in_1 ? 8'h60 : _GEN_303; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_305 = 8'h31 == io_in_1 ? 8'h62 : _GEN_304; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_306 = 8'h32 == io_in_1 ? 8'h64 : _GEN_305; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_307 = 8'h33 == io_in_1 ? 8'h66 : _GEN_306; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_308 = 8'h34 == io_in_1 ? 8'h68 : _GEN_307; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_309 = 8'h35 == io_in_1 ? 8'h6a : _GEN_308; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_310 = 8'h36 == io_in_1 ? 8'h6c : _GEN_309; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_311 = 8'h37 == io_in_1 ? 8'h6e : _GEN_310; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_312 = 8'h38 == io_in_1 ? 8'h70 : _GEN_311; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_313 = 8'h39 == io_in_1 ? 8'h72 : _GEN_312; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_314 = 8'h3a == io_in_1 ? 8'h74 : _GEN_313; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_315 = 8'h3b == io_in_1 ? 8'h76 : _GEN_314; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_316 = 8'h3c == io_in_1 ? 8'h78 : _GEN_315; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_317 = 8'h3d == io_in_1 ? 8'h7a : _GEN_316; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_318 = 8'h3e == io_in_1 ? 8'h7c : _GEN_317; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_319 = 8'h3f == io_in_1 ? 8'h7e : _GEN_318; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_320 = 8'h40 == io_in_1 ? 8'h80 : _GEN_319; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_321 = 8'h41 == io_in_1 ? 8'h82 : _GEN_320; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_322 = 8'h42 == io_in_1 ? 8'h84 : _GEN_321; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_323 = 8'h43 == io_in_1 ? 8'h86 : _GEN_322; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_324 = 8'h44 == io_in_1 ? 8'h88 : _GEN_323; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_325 = 8'h45 == io_in_1 ? 8'h8a : _GEN_324; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_326 = 8'h46 == io_in_1 ? 8'h8c : _GEN_325; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_327 = 8'h47 == io_in_1 ? 8'h8e : _GEN_326; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_328 = 8'h48 == io_in_1 ? 8'h90 : _GEN_327; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_329 = 8'h49 == io_in_1 ? 8'h92 : _GEN_328; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_330 = 8'h4a == io_in_1 ? 8'h94 : _GEN_329; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_331 = 8'h4b == io_in_1 ? 8'h96 : _GEN_330; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_332 = 8'h4c == io_in_1 ? 8'h98 : _GEN_331; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_333 = 8'h4d == io_in_1 ? 8'h9a : _GEN_332; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_334 = 8'h4e == io_in_1 ? 8'h9c : _GEN_333; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_335 = 8'h4f == io_in_1 ? 8'h9e : _GEN_334; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_336 = 8'h50 == io_in_1 ? 8'ha0 : _GEN_335; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_337 = 8'h51 == io_in_1 ? 8'ha2 : _GEN_336; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_338 = 8'h52 == io_in_1 ? 8'ha4 : _GEN_337; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_339 = 8'h53 == io_in_1 ? 8'ha6 : _GEN_338; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_340 = 8'h54 == io_in_1 ? 8'ha8 : _GEN_339; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_341 = 8'h55 == io_in_1 ? 8'haa : _GEN_340; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_342 = 8'h56 == io_in_1 ? 8'hac : _GEN_341; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_343 = 8'h57 == io_in_1 ? 8'hae : _GEN_342; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_344 = 8'h58 == io_in_1 ? 8'hb0 : _GEN_343; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_345 = 8'h59 == io_in_1 ? 8'hb2 : _GEN_344; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_346 = 8'h5a == io_in_1 ? 8'hb4 : _GEN_345; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_347 = 8'h5b == io_in_1 ? 8'hb6 : _GEN_346; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_348 = 8'h5c == io_in_1 ? 8'hb8 : _GEN_347; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_349 = 8'h5d == io_in_1 ? 8'hba : _GEN_348; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_350 = 8'h5e == io_in_1 ? 8'hbc : _GEN_349; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_351 = 8'h5f == io_in_1 ? 8'hbe : _GEN_350; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_352 = 8'h60 == io_in_1 ? 8'hc0 : _GEN_351; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_353 = 8'h61 == io_in_1 ? 8'hc2 : _GEN_352; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_354 = 8'h62 == io_in_1 ? 8'hc4 : _GEN_353; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_355 = 8'h63 == io_in_1 ? 8'hc6 : _GEN_354; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_356 = 8'h64 == io_in_1 ? 8'hc8 : _GEN_355; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_357 = 8'h65 == io_in_1 ? 8'hca : _GEN_356; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_358 = 8'h66 == io_in_1 ? 8'hcc : _GEN_357; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_359 = 8'h67 == io_in_1 ? 8'hce : _GEN_358; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_360 = 8'h68 == io_in_1 ? 8'hd0 : _GEN_359; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_361 = 8'h69 == io_in_1 ? 8'hd2 : _GEN_360; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_362 = 8'h6a == io_in_1 ? 8'hd4 : _GEN_361; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_363 = 8'h6b == io_in_1 ? 8'hd6 : _GEN_362; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_364 = 8'h6c == io_in_1 ? 8'hd8 : _GEN_363; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_365 = 8'h6d == io_in_1 ? 8'hda : _GEN_364; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_366 = 8'h6e == io_in_1 ? 8'hdc : _GEN_365; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_367 = 8'h6f == io_in_1 ? 8'hde : _GEN_366; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_368 = 8'h70 == io_in_1 ? 8'he0 : _GEN_367; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_369 = 8'h71 == io_in_1 ? 8'he2 : _GEN_368; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_370 = 8'h72 == io_in_1 ? 8'he4 : _GEN_369; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_371 = 8'h73 == io_in_1 ? 8'he6 : _GEN_370; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_372 = 8'h74 == io_in_1 ? 8'he8 : _GEN_371; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_373 = 8'h75 == io_in_1 ? 8'hea : _GEN_372; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_374 = 8'h76 == io_in_1 ? 8'hec : _GEN_373; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_375 = 8'h77 == io_in_1 ? 8'hee : _GEN_374; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_376 = 8'h78 == io_in_1 ? 8'hf0 : _GEN_375; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_377 = 8'h79 == io_in_1 ? 8'hf2 : _GEN_376; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_378 = 8'h7a == io_in_1 ? 8'hf4 : _GEN_377; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_379 = 8'h7b == io_in_1 ? 8'hf6 : _GEN_378; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_380 = 8'h7c == io_in_1 ? 8'hf8 : _GEN_379; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_381 = 8'h7d == io_in_1 ? 8'hfa : _GEN_380; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_382 = 8'h7e == io_in_1 ? 8'hfc : _GEN_381; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_383 = 8'h7f == io_in_1 ? 8'hfe : _GEN_382; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_384 = 8'h80 == io_in_1 ? 8'h1b : _GEN_383; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_385 = 8'h81 == io_in_1 ? 8'h19 : _GEN_384; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_386 = 8'h82 == io_in_1 ? 8'h1f : _GEN_385; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_387 = 8'h83 == io_in_1 ? 8'h1d : _GEN_386; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_388 = 8'h84 == io_in_1 ? 8'h13 : _GEN_387; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_389 = 8'h85 == io_in_1 ? 8'h11 : _GEN_388; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_390 = 8'h86 == io_in_1 ? 8'h17 : _GEN_389; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_391 = 8'h87 == io_in_1 ? 8'h15 : _GEN_390; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_392 = 8'h88 == io_in_1 ? 8'hb : _GEN_391; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_393 = 8'h89 == io_in_1 ? 8'h9 : _GEN_392; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_394 = 8'h8a == io_in_1 ? 8'hf : _GEN_393; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_395 = 8'h8b == io_in_1 ? 8'hd : _GEN_394; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_396 = 8'h8c == io_in_1 ? 8'h3 : _GEN_395; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_397 = 8'h8d == io_in_1 ? 8'h1 : _GEN_396; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_398 = 8'h8e == io_in_1 ? 8'h7 : _GEN_397; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_399 = 8'h8f == io_in_1 ? 8'h5 : _GEN_398; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_400 = 8'h90 == io_in_1 ? 8'h3b : _GEN_399; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_401 = 8'h91 == io_in_1 ? 8'h39 : _GEN_400; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_402 = 8'h92 == io_in_1 ? 8'h3f : _GEN_401; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_403 = 8'h93 == io_in_1 ? 8'h3d : _GEN_402; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_404 = 8'h94 == io_in_1 ? 8'h33 : _GEN_403; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_405 = 8'h95 == io_in_1 ? 8'h31 : _GEN_404; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_406 = 8'h96 == io_in_1 ? 8'h37 : _GEN_405; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_407 = 8'h97 == io_in_1 ? 8'h35 : _GEN_406; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_408 = 8'h98 == io_in_1 ? 8'h2b : _GEN_407; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_409 = 8'h99 == io_in_1 ? 8'h29 : _GEN_408; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_410 = 8'h9a == io_in_1 ? 8'h2f : _GEN_409; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_411 = 8'h9b == io_in_1 ? 8'h2d : _GEN_410; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_412 = 8'h9c == io_in_1 ? 8'h23 : _GEN_411; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_413 = 8'h9d == io_in_1 ? 8'h21 : _GEN_412; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_414 = 8'h9e == io_in_1 ? 8'h27 : _GEN_413; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_415 = 8'h9f == io_in_1 ? 8'h25 : _GEN_414; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_416 = 8'ha0 == io_in_1 ? 8'h5b : _GEN_415; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_417 = 8'ha1 == io_in_1 ? 8'h59 : _GEN_416; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_418 = 8'ha2 == io_in_1 ? 8'h5f : _GEN_417; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_419 = 8'ha3 == io_in_1 ? 8'h5d : _GEN_418; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_420 = 8'ha4 == io_in_1 ? 8'h53 : _GEN_419; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_421 = 8'ha5 == io_in_1 ? 8'h51 : _GEN_420; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_422 = 8'ha6 == io_in_1 ? 8'h57 : _GEN_421; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_423 = 8'ha7 == io_in_1 ? 8'h55 : _GEN_422; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_424 = 8'ha8 == io_in_1 ? 8'h4b : _GEN_423; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_425 = 8'ha9 == io_in_1 ? 8'h49 : _GEN_424; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_426 = 8'haa == io_in_1 ? 8'h4f : _GEN_425; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_427 = 8'hab == io_in_1 ? 8'h4d : _GEN_426; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_428 = 8'hac == io_in_1 ? 8'h43 : _GEN_427; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_429 = 8'had == io_in_1 ? 8'h41 : _GEN_428; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_430 = 8'hae == io_in_1 ? 8'h47 : _GEN_429; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_431 = 8'haf == io_in_1 ? 8'h45 : _GEN_430; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_432 = 8'hb0 == io_in_1 ? 8'h7b : _GEN_431; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_433 = 8'hb1 == io_in_1 ? 8'h79 : _GEN_432; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_434 = 8'hb2 == io_in_1 ? 8'h7f : _GEN_433; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_435 = 8'hb3 == io_in_1 ? 8'h7d : _GEN_434; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_436 = 8'hb4 == io_in_1 ? 8'h73 : _GEN_435; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_437 = 8'hb5 == io_in_1 ? 8'h71 : _GEN_436; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_438 = 8'hb6 == io_in_1 ? 8'h77 : _GEN_437; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_439 = 8'hb7 == io_in_1 ? 8'h75 : _GEN_438; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_440 = 8'hb8 == io_in_1 ? 8'h6b : _GEN_439; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_441 = 8'hb9 == io_in_1 ? 8'h69 : _GEN_440; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_442 = 8'hba == io_in_1 ? 8'h6f : _GEN_441; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_443 = 8'hbb == io_in_1 ? 8'h6d : _GEN_442; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_444 = 8'hbc == io_in_1 ? 8'h63 : _GEN_443; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_445 = 8'hbd == io_in_1 ? 8'h61 : _GEN_444; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_446 = 8'hbe == io_in_1 ? 8'h67 : _GEN_445; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_447 = 8'hbf == io_in_1 ? 8'h65 : _GEN_446; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_448 = 8'hc0 == io_in_1 ? 8'h9b : _GEN_447; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_449 = 8'hc1 == io_in_1 ? 8'h99 : _GEN_448; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_450 = 8'hc2 == io_in_1 ? 8'h9f : _GEN_449; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_451 = 8'hc3 == io_in_1 ? 8'h9d : _GEN_450; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_452 = 8'hc4 == io_in_1 ? 8'h93 : _GEN_451; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_453 = 8'hc5 == io_in_1 ? 8'h91 : _GEN_452; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_454 = 8'hc6 == io_in_1 ? 8'h97 : _GEN_453; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_455 = 8'hc7 == io_in_1 ? 8'h95 : _GEN_454; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_456 = 8'hc8 == io_in_1 ? 8'h8b : _GEN_455; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_457 = 8'hc9 == io_in_1 ? 8'h89 : _GEN_456; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_458 = 8'hca == io_in_1 ? 8'h8f : _GEN_457; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_459 = 8'hcb == io_in_1 ? 8'h8d : _GEN_458; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_460 = 8'hcc == io_in_1 ? 8'h83 : _GEN_459; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_461 = 8'hcd == io_in_1 ? 8'h81 : _GEN_460; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_462 = 8'hce == io_in_1 ? 8'h87 : _GEN_461; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_463 = 8'hcf == io_in_1 ? 8'h85 : _GEN_462; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_464 = 8'hd0 == io_in_1 ? 8'hbb : _GEN_463; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_465 = 8'hd1 == io_in_1 ? 8'hb9 : _GEN_464; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_466 = 8'hd2 == io_in_1 ? 8'hbf : _GEN_465; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_467 = 8'hd3 == io_in_1 ? 8'hbd : _GEN_466; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_468 = 8'hd4 == io_in_1 ? 8'hb3 : _GEN_467; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_469 = 8'hd5 == io_in_1 ? 8'hb1 : _GEN_468; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_470 = 8'hd6 == io_in_1 ? 8'hb7 : _GEN_469; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_471 = 8'hd7 == io_in_1 ? 8'hb5 : _GEN_470; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_472 = 8'hd8 == io_in_1 ? 8'hab : _GEN_471; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_473 = 8'hd9 == io_in_1 ? 8'ha9 : _GEN_472; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_474 = 8'hda == io_in_1 ? 8'haf : _GEN_473; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_475 = 8'hdb == io_in_1 ? 8'had : _GEN_474; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_476 = 8'hdc == io_in_1 ? 8'ha3 : _GEN_475; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_477 = 8'hdd == io_in_1 ? 8'ha1 : _GEN_476; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_478 = 8'hde == io_in_1 ? 8'ha7 : _GEN_477; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_479 = 8'hdf == io_in_1 ? 8'ha5 : _GEN_478; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_480 = 8'he0 == io_in_1 ? 8'hdb : _GEN_479; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_481 = 8'he1 == io_in_1 ? 8'hd9 : _GEN_480; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_482 = 8'he2 == io_in_1 ? 8'hdf : _GEN_481; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_483 = 8'he3 == io_in_1 ? 8'hdd : _GEN_482; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_484 = 8'he4 == io_in_1 ? 8'hd3 : _GEN_483; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_485 = 8'he5 == io_in_1 ? 8'hd1 : _GEN_484; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_486 = 8'he6 == io_in_1 ? 8'hd7 : _GEN_485; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_487 = 8'he7 == io_in_1 ? 8'hd5 : _GEN_486; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_488 = 8'he8 == io_in_1 ? 8'hcb : _GEN_487; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_489 = 8'he9 == io_in_1 ? 8'hc9 : _GEN_488; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_490 = 8'hea == io_in_1 ? 8'hcf : _GEN_489; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_491 = 8'heb == io_in_1 ? 8'hcd : _GEN_490; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_492 = 8'hec == io_in_1 ? 8'hc3 : _GEN_491; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_493 = 8'hed == io_in_1 ? 8'hc1 : _GEN_492; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_494 = 8'hee == io_in_1 ? 8'hc7 : _GEN_493; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_495 = 8'hef == io_in_1 ? 8'hc5 : _GEN_494; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_496 = 8'hf0 == io_in_1 ? 8'hfb : _GEN_495; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_497 = 8'hf1 == io_in_1 ? 8'hf9 : _GEN_496; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_498 = 8'hf2 == io_in_1 ? 8'hff : _GEN_497; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_499 = 8'hf3 == io_in_1 ? 8'hfd : _GEN_498; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_500 = 8'hf4 == io_in_1 ? 8'hf3 : _GEN_499; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_501 = 8'hf5 == io_in_1 ? 8'hf1 : _GEN_500; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_502 = 8'hf6 == io_in_1 ? 8'hf7 : _GEN_501; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_503 = 8'hf7 == io_in_1 ? 8'hf5 : _GEN_502; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_504 = 8'hf8 == io_in_1 ? 8'heb : _GEN_503; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_505 = 8'hf9 == io_in_1 ? 8'he9 : _GEN_504; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_506 = 8'hfa == io_in_1 ? 8'hef : _GEN_505; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_507 = 8'hfb == io_in_1 ? 8'hed : _GEN_506; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_508 = 8'hfc == io_in_1 ? 8'he3 : _GEN_507; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_509 = 8'hfd == io_in_1 ? 8'he1 : _GEN_508; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_510 = 8'hfe == io_in_1 ? 8'he7 : _GEN_509; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _GEN_511 = 8'hff == io_in_1 ? 8'he5 : _GEN_510; // @[AES_PipelinedElasticBuffer.scala 328:31 AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _T = _GEN_255 ^ _GEN_511; // @[AES_PipelinedElasticBuffer.scala 328:31]
  wire [7:0] _T_1 = _T ^ io_in_1; // @[AES_PipelinedElasticBuffer.scala 328:48]
  wire [7:0] _T_2 = _T_1 ^ io_in_2; // @[AES_PipelinedElasticBuffer.scala 328:59]
  wire [7:0] _T_4 = io_in_0 ^ _GEN_511; // @[AES_PipelinedElasticBuffer.scala 329:25]
  wire [7:0] _GEN_513 = 8'h1 == io_in_2 ? 8'h2 : 8'h0; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_514 = 8'h2 == io_in_2 ? 8'h4 : _GEN_513; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_515 = 8'h3 == io_in_2 ? 8'h6 : _GEN_514; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_516 = 8'h4 == io_in_2 ? 8'h8 : _GEN_515; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_517 = 8'h5 == io_in_2 ? 8'ha : _GEN_516; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_518 = 8'h6 == io_in_2 ? 8'hc : _GEN_517; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_519 = 8'h7 == io_in_2 ? 8'he : _GEN_518; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_520 = 8'h8 == io_in_2 ? 8'h10 : _GEN_519; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_521 = 8'h9 == io_in_2 ? 8'h12 : _GEN_520; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_522 = 8'ha == io_in_2 ? 8'h14 : _GEN_521; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_523 = 8'hb == io_in_2 ? 8'h16 : _GEN_522; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_524 = 8'hc == io_in_2 ? 8'h18 : _GEN_523; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_525 = 8'hd == io_in_2 ? 8'h1a : _GEN_524; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_526 = 8'he == io_in_2 ? 8'h1c : _GEN_525; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_527 = 8'hf == io_in_2 ? 8'h1e : _GEN_526; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_528 = 8'h10 == io_in_2 ? 8'h20 : _GEN_527; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_529 = 8'h11 == io_in_2 ? 8'h22 : _GEN_528; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_530 = 8'h12 == io_in_2 ? 8'h24 : _GEN_529; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_531 = 8'h13 == io_in_2 ? 8'h26 : _GEN_530; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_532 = 8'h14 == io_in_2 ? 8'h28 : _GEN_531; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_533 = 8'h15 == io_in_2 ? 8'h2a : _GEN_532; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_534 = 8'h16 == io_in_2 ? 8'h2c : _GEN_533; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_535 = 8'h17 == io_in_2 ? 8'h2e : _GEN_534; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_536 = 8'h18 == io_in_2 ? 8'h30 : _GEN_535; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_537 = 8'h19 == io_in_2 ? 8'h32 : _GEN_536; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_538 = 8'h1a == io_in_2 ? 8'h34 : _GEN_537; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_539 = 8'h1b == io_in_2 ? 8'h36 : _GEN_538; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_540 = 8'h1c == io_in_2 ? 8'h38 : _GEN_539; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_541 = 8'h1d == io_in_2 ? 8'h3a : _GEN_540; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_542 = 8'h1e == io_in_2 ? 8'h3c : _GEN_541; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_543 = 8'h1f == io_in_2 ? 8'h3e : _GEN_542; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_544 = 8'h20 == io_in_2 ? 8'h40 : _GEN_543; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_545 = 8'h21 == io_in_2 ? 8'h42 : _GEN_544; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_546 = 8'h22 == io_in_2 ? 8'h44 : _GEN_545; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_547 = 8'h23 == io_in_2 ? 8'h46 : _GEN_546; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_548 = 8'h24 == io_in_2 ? 8'h48 : _GEN_547; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_549 = 8'h25 == io_in_2 ? 8'h4a : _GEN_548; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_550 = 8'h26 == io_in_2 ? 8'h4c : _GEN_549; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_551 = 8'h27 == io_in_2 ? 8'h4e : _GEN_550; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_552 = 8'h28 == io_in_2 ? 8'h50 : _GEN_551; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_553 = 8'h29 == io_in_2 ? 8'h52 : _GEN_552; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_554 = 8'h2a == io_in_2 ? 8'h54 : _GEN_553; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_555 = 8'h2b == io_in_2 ? 8'h56 : _GEN_554; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_556 = 8'h2c == io_in_2 ? 8'h58 : _GEN_555; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_557 = 8'h2d == io_in_2 ? 8'h5a : _GEN_556; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_558 = 8'h2e == io_in_2 ? 8'h5c : _GEN_557; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_559 = 8'h2f == io_in_2 ? 8'h5e : _GEN_558; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_560 = 8'h30 == io_in_2 ? 8'h60 : _GEN_559; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_561 = 8'h31 == io_in_2 ? 8'h62 : _GEN_560; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_562 = 8'h32 == io_in_2 ? 8'h64 : _GEN_561; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_563 = 8'h33 == io_in_2 ? 8'h66 : _GEN_562; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_564 = 8'h34 == io_in_2 ? 8'h68 : _GEN_563; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_565 = 8'h35 == io_in_2 ? 8'h6a : _GEN_564; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_566 = 8'h36 == io_in_2 ? 8'h6c : _GEN_565; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_567 = 8'h37 == io_in_2 ? 8'h6e : _GEN_566; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_568 = 8'h38 == io_in_2 ? 8'h70 : _GEN_567; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_569 = 8'h39 == io_in_2 ? 8'h72 : _GEN_568; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_570 = 8'h3a == io_in_2 ? 8'h74 : _GEN_569; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_571 = 8'h3b == io_in_2 ? 8'h76 : _GEN_570; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_572 = 8'h3c == io_in_2 ? 8'h78 : _GEN_571; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_573 = 8'h3d == io_in_2 ? 8'h7a : _GEN_572; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_574 = 8'h3e == io_in_2 ? 8'h7c : _GEN_573; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_575 = 8'h3f == io_in_2 ? 8'h7e : _GEN_574; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_576 = 8'h40 == io_in_2 ? 8'h80 : _GEN_575; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_577 = 8'h41 == io_in_2 ? 8'h82 : _GEN_576; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_578 = 8'h42 == io_in_2 ? 8'h84 : _GEN_577; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_579 = 8'h43 == io_in_2 ? 8'h86 : _GEN_578; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_580 = 8'h44 == io_in_2 ? 8'h88 : _GEN_579; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_581 = 8'h45 == io_in_2 ? 8'h8a : _GEN_580; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_582 = 8'h46 == io_in_2 ? 8'h8c : _GEN_581; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_583 = 8'h47 == io_in_2 ? 8'h8e : _GEN_582; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_584 = 8'h48 == io_in_2 ? 8'h90 : _GEN_583; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_585 = 8'h49 == io_in_2 ? 8'h92 : _GEN_584; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_586 = 8'h4a == io_in_2 ? 8'h94 : _GEN_585; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_587 = 8'h4b == io_in_2 ? 8'h96 : _GEN_586; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_588 = 8'h4c == io_in_2 ? 8'h98 : _GEN_587; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_589 = 8'h4d == io_in_2 ? 8'h9a : _GEN_588; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_590 = 8'h4e == io_in_2 ? 8'h9c : _GEN_589; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_591 = 8'h4f == io_in_2 ? 8'h9e : _GEN_590; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_592 = 8'h50 == io_in_2 ? 8'ha0 : _GEN_591; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_593 = 8'h51 == io_in_2 ? 8'ha2 : _GEN_592; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_594 = 8'h52 == io_in_2 ? 8'ha4 : _GEN_593; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_595 = 8'h53 == io_in_2 ? 8'ha6 : _GEN_594; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_596 = 8'h54 == io_in_2 ? 8'ha8 : _GEN_595; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_597 = 8'h55 == io_in_2 ? 8'haa : _GEN_596; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_598 = 8'h56 == io_in_2 ? 8'hac : _GEN_597; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_599 = 8'h57 == io_in_2 ? 8'hae : _GEN_598; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_600 = 8'h58 == io_in_2 ? 8'hb0 : _GEN_599; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_601 = 8'h59 == io_in_2 ? 8'hb2 : _GEN_600; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_602 = 8'h5a == io_in_2 ? 8'hb4 : _GEN_601; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_603 = 8'h5b == io_in_2 ? 8'hb6 : _GEN_602; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_604 = 8'h5c == io_in_2 ? 8'hb8 : _GEN_603; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_605 = 8'h5d == io_in_2 ? 8'hba : _GEN_604; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_606 = 8'h5e == io_in_2 ? 8'hbc : _GEN_605; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_607 = 8'h5f == io_in_2 ? 8'hbe : _GEN_606; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_608 = 8'h60 == io_in_2 ? 8'hc0 : _GEN_607; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_609 = 8'h61 == io_in_2 ? 8'hc2 : _GEN_608; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_610 = 8'h62 == io_in_2 ? 8'hc4 : _GEN_609; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_611 = 8'h63 == io_in_2 ? 8'hc6 : _GEN_610; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_612 = 8'h64 == io_in_2 ? 8'hc8 : _GEN_611; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_613 = 8'h65 == io_in_2 ? 8'hca : _GEN_612; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_614 = 8'h66 == io_in_2 ? 8'hcc : _GEN_613; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_615 = 8'h67 == io_in_2 ? 8'hce : _GEN_614; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_616 = 8'h68 == io_in_2 ? 8'hd0 : _GEN_615; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_617 = 8'h69 == io_in_2 ? 8'hd2 : _GEN_616; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_618 = 8'h6a == io_in_2 ? 8'hd4 : _GEN_617; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_619 = 8'h6b == io_in_2 ? 8'hd6 : _GEN_618; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_620 = 8'h6c == io_in_2 ? 8'hd8 : _GEN_619; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_621 = 8'h6d == io_in_2 ? 8'hda : _GEN_620; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_622 = 8'h6e == io_in_2 ? 8'hdc : _GEN_621; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_623 = 8'h6f == io_in_2 ? 8'hde : _GEN_622; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_624 = 8'h70 == io_in_2 ? 8'he0 : _GEN_623; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_625 = 8'h71 == io_in_2 ? 8'he2 : _GEN_624; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_626 = 8'h72 == io_in_2 ? 8'he4 : _GEN_625; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_627 = 8'h73 == io_in_2 ? 8'he6 : _GEN_626; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_628 = 8'h74 == io_in_2 ? 8'he8 : _GEN_627; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_629 = 8'h75 == io_in_2 ? 8'hea : _GEN_628; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_630 = 8'h76 == io_in_2 ? 8'hec : _GEN_629; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_631 = 8'h77 == io_in_2 ? 8'hee : _GEN_630; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_632 = 8'h78 == io_in_2 ? 8'hf0 : _GEN_631; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_633 = 8'h79 == io_in_2 ? 8'hf2 : _GEN_632; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_634 = 8'h7a == io_in_2 ? 8'hf4 : _GEN_633; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_635 = 8'h7b == io_in_2 ? 8'hf6 : _GEN_634; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_636 = 8'h7c == io_in_2 ? 8'hf8 : _GEN_635; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_637 = 8'h7d == io_in_2 ? 8'hfa : _GEN_636; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_638 = 8'h7e == io_in_2 ? 8'hfc : _GEN_637; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_639 = 8'h7f == io_in_2 ? 8'hfe : _GEN_638; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_640 = 8'h80 == io_in_2 ? 8'h1b : _GEN_639; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_641 = 8'h81 == io_in_2 ? 8'h19 : _GEN_640; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_642 = 8'h82 == io_in_2 ? 8'h1f : _GEN_641; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_643 = 8'h83 == io_in_2 ? 8'h1d : _GEN_642; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_644 = 8'h84 == io_in_2 ? 8'h13 : _GEN_643; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_645 = 8'h85 == io_in_2 ? 8'h11 : _GEN_644; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_646 = 8'h86 == io_in_2 ? 8'h17 : _GEN_645; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_647 = 8'h87 == io_in_2 ? 8'h15 : _GEN_646; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_648 = 8'h88 == io_in_2 ? 8'hb : _GEN_647; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_649 = 8'h89 == io_in_2 ? 8'h9 : _GEN_648; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_650 = 8'h8a == io_in_2 ? 8'hf : _GEN_649; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_651 = 8'h8b == io_in_2 ? 8'hd : _GEN_650; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_652 = 8'h8c == io_in_2 ? 8'h3 : _GEN_651; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_653 = 8'h8d == io_in_2 ? 8'h1 : _GEN_652; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_654 = 8'h8e == io_in_2 ? 8'h7 : _GEN_653; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_655 = 8'h8f == io_in_2 ? 8'h5 : _GEN_654; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_656 = 8'h90 == io_in_2 ? 8'h3b : _GEN_655; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_657 = 8'h91 == io_in_2 ? 8'h39 : _GEN_656; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_658 = 8'h92 == io_in_2 ? 8'h3f : _GEN_657; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_659 = 8'h93 == io_in_2 ? 8'h3d : _GEN_658; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_660 = 8'h94 == io_in_2 ? 8'h33 : _GEN_659; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_661 = 8'h95 == io_in_2 ? 8'h31 : _GEN_660; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_662 = 8'h96 == io_in_2 ? 8'h37 : _GEN_661; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_663 = 8'h97 == io_in_2 ? 8'h35 : _GEN_662; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_664 = 8'h98 == io_in_2 ? 8'h2b : _GEN_663; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_665 = 8'h99 == io_in_2 ? 8'h29 : _GEN_664; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_666 = 8'h9a == io_in_2 ? 8'h2f : _GEN_665; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_667 = 8'h9b == io_in_2 ? 8'h2d : _GEN_666; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_668 = 8'h9c == io_in_2 ? 8'h23 : _GEN_667; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_669 = 8'h9d == io_in_2 ? 8'h21 : _GEN_668; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_670 = 8'h9e == io_in_2 ? 8'h27 : _GEN_669; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_671 = 8'h9f == io_in_2 ? 8'h25 : _GEN_670; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_672 = 8'ha0 == io_in_2 ? 8'h5b : _GEN_671; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_673 = 8'ha1 == io_in_2 ? 8'h59 : _GEN_672; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_674 = 8'ha2 == io_in_2 ? 8'h5f : _GEN_673; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_675 = 8'ha3 == io_in_2 ? 8'h5d : _GEN_674; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_676 = 8'ha4 == io_in_2 ? 8'h53 : _GEN_675; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_677 = 8'ha5 == io_in_2 ? 8'h51 : _GEN_676; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_678 = 8'ha6 == io_in_2 ? 8'h57 : _GEN_677; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_679 = 8'ha7 == io_in_2 ? 8'h55 : _GEN_678; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_680 = 8'ha8 == io_in_2 ? 8'h4b : _GEN_679; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_681 = 8'ha9 == io_in_2 ? 8'h49 : _GEN_680; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_682 = 8'haa == io_in_2 ? 8'h4f : _GEN_681; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_683 = 8'hab == io_in_2 ? 8'h4d : _GEN_682; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_684 = 8'hac == io_in_2 ? 8'h43 : _GEN_683; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_685 = 8'had == io_in_2 ? 8'h41 : _GEN_684; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_686 = 8'hae == io_in_2 ? 8'h47 : _GEN_685; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_687 = 8'haf == io_in_2 ? 8'h45 : _GEN_686; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_688 = 8'hb0 == io_in_2 ? 8'h7b : _GEN_687; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_689 = 8'hb1 == io_in_2 ? 8'h79 : _GEN_688; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_690 = 8'hb2 == io_in_2 ? 8'h7f : _GEN_689; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_691 = 8'hb3 == io_in_2 ? 8'h7d : _GEN_690; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_692 = 8'hb4 == io_in_2 ? 8'h73 : _GEN_691; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_693 = 8'hb5 == io_in_2 ? 8'h71 : _GEN_692; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_694 = 8'hb6 == io_in_2 ? 8'h77 : _GEN_693; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_695 = 8'hb7 == io_in_2 ? 8'h75 : _GEN_694; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_696 = 8'hb8 == io_in_2 ? 8'h6b : _GEN_695; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_697 = 8'hb9 == io_in_2 ? 8'h69 : _GEN_696; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_698 = 8'hba == io_in_2 ? 8'h6f : _GEN_697; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_699 = 8'hbb == io_in_2 ? 8'h6d : _GEN_698; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_700 = 8'hbc == io_in_2 ? 8'h63 : _GEN_699; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_701 = 8'hbd == io_in_2 ? 8'h61 : _GEN_700; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_702 = 8'hbe == io_in_2 ? 8'h67 : _GEN_701; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_703 = 8'hbf == io_in_2 ? 8'h65 : _GEN_702; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_704 = 8'hc0 == io_in_2 ? 8'h9b : _GEN_703; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_705 = 8'hc1 == io_in_2 ? 8'h99 : _GEN_704; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_706 = 8'hc2 == io_in_2 ? 8'h9f : _GEN_705; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_707 = 8'hc3 == io_in_2 ? 8'h9d : _GEN_706; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_708 = 8'hc4 == io_in_2 ? 8'h93 : _GEN_707; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_709 = 8'hc5 == io_in_2 ? 8'h91 : _GEN_708; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_710 = 8'hc6 == io_in_2 ? 8'h97 : _GEN_709; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_711 = 8'hc7 == io_in_2 ? 8'h95 : _GEN_710; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_712 = 8'hc8 == io_in_2 ? 8'h8b : _GEN_711; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_713 = 8'hc9 == io_in_2 ? 8'h89 : _GEN_712; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_714 = 8'hca == io_in_2 ? 8'h8f : _GEN_713; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_715 = 8'hcb == io_in_2 ? 8'h8d : _GEN_714; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_716 = 8'hcc == io_in_2 ? 8'h83 : _GEN_715; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_717 = 8'hcd == io_in_2 ? 8'h81 : _GEN_716; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_718 = 8'hce == io_in_2 ? 8'h87 : _GEN_717; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_719 = 8'hcf == io_in_2 ? 8'h85 : _GEN_718; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_720 = 8'hd0 == io_in_2 ? 8'hbb : _GEN_719; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_721 = 8'hd1 == io_in_2 ? 8'hb9 : _GEN_720; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_722 = 8'hd2 == io_in_2 ? 8'hbf : _GEN_721; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_723 = 8'hd3 == io_in_2 ? 8'hbd : _GEN_722; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_724 = 8'hd4 == io_in_2 ? 8'hb3 : _GEN_723; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_725 = 8'hd5 == io_in_2 ? 8'hb1 : _GEN_724; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_726 = 8'hd6 == io_in_2 ? 8'hb7 : _GEN_725; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_727 = 8'hd7 == io_in_2 ? 8'hb5 : _GEN_726; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_728 = 8'hd8 == io_in_2 ? 8'hab : _GEN_727; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_729 = 8'hd9 == io_in_2 ? 8'ha9 : _GEN_728; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_730 = 8'hda == io_in_2 ? 8'haf : _GEN_729; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_731 = 8'hdb == io_in_2 ? 8'had : _GEN_730; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_732 = 8'hdc == io_in_2 ? 8'ha3 : _GEN_731; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_733 = 8'hdd == io_in_2 ? 8'ha1 : _GEN_732; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_734 = 8'hde == io_in_2 ? 8'ha7 : _GEN_733; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_735 = 8'hdf == io_in_2 ? 8'ha5 : _GEN_734; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_736 = 8'he0 == io_in_2 ? 8'hdb : _GEN_735; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_737 = 8'he1 == io_in_2 ? 8'hd9 : _GEN_736; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_738 = 8'he2 == io_in_2 ? 8'hdf : _GEN_737; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_739 = 8'he3 == io_in_2 ? 8'hdd : _GEN_738; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_740 = 8'he4 == io_in_2 ? 8'hd3 : _GEN_739; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_741 = 8'he5 == io_in_2 ? 8'hd1 : _GEN_740; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_742 = 8'he6 == io_in_2 ? 8'hd7 : _GEN_741; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_743 = 8'he7 == io_in_2 ? 8'hd5 : _GEN_742; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_744 = 8'he8 == io_in_2 ? 8'hcb : _GEN_743; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_745 = 8'he9 == io_in_2 ? 8'hc9 : _GEN_744; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_746 = 8'hea == io_in_2 ? 8'hcf : _GEN_745; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_747 = 8'heb == io_in_2 ? 8'hcd : _GEN_746; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_748 = 8'hec == io_in_2 ? 8'hc3 : _GEN_747; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_749 = 8'hed == io_in_2 ? 8'hc1 : _GEN_748; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_750 = 8'hee == io_in_2 ? 8'hc7 : _GEN_749; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_751 = 8'hef == io_in_2 ? 8'hc5 : _GEN_750; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_752 = 8'hf0 == io_in_2 ? 8'hfb : _GEN_751; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_753 = 8'hf1 == io_in_2 ? 8'hf9 : _GEN_752; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_754 = 8'hf2 == io_in_2 ? 8'hff : _GEN_753; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_755 = 8'hf3 == io_in_2 ? 8'hfd : _GEN_754; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_756 = 8'hf4 == io_in_2 ? 8'hf3 : _GEN_755; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_757 = 8'hf5 == io_in_2 ? 8'hf1 : _GEN_756; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_758 = 8'hf6 == io_in_2 ? 8'hf7 : _GEN_757; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_759 = 8'hf7 == io_in_2 ? 8'hf5 : _GEN_758; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_760 = 8'hf8 == io_in_2 ? 8'heb : _GEN_759; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_761 = 8'hf9 == io_in_2 ? 8'he9 : _GEN_760; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_762 = 8'hfa == io_in_2 ? 8'hef : _GEN_761; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_763 = 8'hfb == io_in_2 ? 8'hed : _GEN_762; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_764 = 8'hfc == io_in_2 ? 8'he3 : _GEN_763; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_765 = 8'hfd == io_in_2 ? 8'he1 : _GEN_764; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_766 = 8'hfe == io_in_2 ? 8'he7 : _GEN_765; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _GEN_767 = 8'hff == io_in_2 ? 8'he5 : _GEN_766; // @[AES_PipelinedElasticBuffer.scala 329:42 AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _T_5 = _T_4 ^ _GEN_767; // @[AES_PipelinedElasticBuffer.scala 329:42]
  wire [7:0] _T_6 = _T_5 ^ io_in_2; // @[AES_PipelinedElasticBuffer.scala 329:59]
  wire [7:0] _T_8 = io_in_0 ^ io_in_1; // @[AES_PipelinedElasticBuffer.scala 330:25]
  wire [7:0] _T_9 = _T_8 ^ _GEN_767; // @[AES_PipelinedElasticBuffer.scala 330:36]
  wire [7:0] _GEN_769 = 8'h1 == io_in_3 ? 8'h2 : 8'h0; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_770 = 8'h2 == io_in_3 ? 8'h4 : _GEN_769; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_771 = 8'h3 == io_in_3 ? 8'h6 : _GEN_770; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_772 = 8'h4 == io_in_3 ? 8'h8 : _GEN_771; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_773 = 8'h5 == io_in_3 ? 8'ha : _GEN_772; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_774 = 8'h6 == io_in_3 ? 8'hc : _GEN_773; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_775 = 8'h7 == io_in_3 ? 8'he : _GEN_774; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_776 = 8'h8 == io_in_3 ? 8'h10 : _GEN_775; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_777 = 8'h9 == io_in_3 ? 8'h12 : _GEN_776; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_778 = 8'ha == io_in_3 ? 8'h14 : _GEN_777; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_779 = 8'hb == io_in_3 ? 8'h16 : _GEN_778; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_780 = 8'hc == io_in_3 ? 8'h18 : _GEN_779; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_781 = 8'hd == io_in_3 ? 8'h1a : _GEN_780; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_782 = 8'he == io_in_3 ? 8'h1c : _GEN_781; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_783 = 8'hf == io_in_3 ? 8'h1e : _GEN_782; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_784 = 8'h10 == io_in_3 ? 8'h20 : _GEN_783; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_785 = 8'h11 == io_in_3 ? 8'h22 : _GEN_784; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_786 = 8'h12 == io_in_3 ? 8'h24 : _GEN_785; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_787 = 8'h13 == io_in_3 ? 8'h26 : _GEN_786; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_788 = 8'h14 == io_in_3 ? 8'h28 : _GEN_787; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_789 = 8'h15 == io_in_3 ? 8'h2a : _GEN_788; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_790 = 8'h16 == io_in_3 ? 8'h2c : _GEN_789; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_791 = 8'h17 == io_in_3 ? 8'h2e : _GEN_790; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_792 = 8'h18 == io_in_3 ? 8'h30 : _GEN_791; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_793 = 8'h19 == io_in_3 ? 8'h32 : _GEN_792; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_794 = 8'h1a == io_in_3 ? 8'h34 : _GEN_793; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_795 = 8'h1b == io_in_3 ? 8'h36 : _GEN_794; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_796 = 8'h1c == io_in_3 ? 8'h38 : _GEN_795; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_797 = 8'h1d == io_in_3 ? 8'h3a : _GEN_796; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_798 = 8'h1e == io_in_3 ? 8'h3c : _GEN_797; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_799 = 8'h1f == io_in_3 ? 8'h3e : _GEN_798; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_800 = 8'h20 == io_in_3 ? 8'h40 : _GEN_799; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_801 = 8'h21 == io_in_3 ? 8'h42 : _GEN_800; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_802 = 8'h22 == io_in_3 ? 8'h44 : _GEN_801; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_803 = 8'h23 == io_in_3 ? 8'h46 : _GEN_802; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_804 = 8'h24 == io_in_3 ? 8'h48 : _GEN_803; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_805 = 8'h25 == io_in_3 ? 8'h4a : _GEN_804; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_806 = 8'h26 == io_in_3 ? 8'h4c : _GEN_805; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_807 = 8'h27 == io_in_3 ? 8'h4e : _GEN_806; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_808 = 8'h28 == io_in_3 ? 8'h50 : _GEN_807; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_809 = 8'h29 == io_in_3 ? 8'h52 : _GEN_808; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_810 = 8'h2a == io_in_3 ? 8'h54 : _GEN_809; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_811 = 8'h2b == io_in_3 ? 8'h56 : _GEN_810; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_812 = 8'h2c == io_in_3 ? 8'h58 : _GEN_811; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_813 = 8'h2d == io_in_3 ? 8'h5a : _GEN_812; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_814 = 8'h2e == io_in_3 ? 8'h5c : _GEN_813; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_815 = 8'h2f == io_in_3 ? 8'h5e : _GEN_814; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_816 = 8'h30 == io_in_3 ? 8'h60 : _GEN_815; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_817 = 8'h31 == io_in_3 ? 8'h62 : _GEN_816; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_818 = 8'h32 == io_in_3 ? 8'h64 : _GEN_817; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_819 = 8'h33 == io_in_3 ? 8'h66 : _GEN_818; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_820 = 8'h34 == io_in_3 ? 8'h68 : _GEN_819; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_821 = 8'h35 == io_in_3 ? 8'h6a : _GEN_820; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_822 = 8'h36 == io_in_3 ? 8'h6c : _GEN_821; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_823 = 8'h37 == io_in_3 ? 8'h6e : _GEN_822; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_824 = 8'h38 == io_in_3 ? 8'h70 : _GEN_823; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_825 = 8'h39 == io_in_3 ? 8'h72 : _GEN_824; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_826 = 8'h3a == io_in_3 ? 8'h74 : _GEN_825; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_827 = 8'h3b == io_in_3 ? 8'h76 : _GEN_826; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_828 = 8'h3c == io_in_3 ? 8'h78 : _GEN_827; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_829 = 8'h3d == io_in_3 ? 8'h7a : _GEN_828; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_830 = 8'h3e == io_in_3 ? 8'h7c : _GEN_829; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_831 = 8'h3f == io_in_3 ? 8'h7e : _GEN_830; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_832 = 8'h40 == io_in_3 ? 8'h80 : _GEN_831; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_833 = 8'h41 == io_in_3 ? 8'h82 : _GEN_832; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_834 = 8'h42 == io_in_3 ? 8'h84 : _GEN_833; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_835 = 8'h43 == io_in_3 ? 8'h86 : _GEN_834; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_836 = 8'h44 == io_in_3 ? 8'h88 : _GEN_835; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_837 = 8'h45 == io_in_3 ? 8'h8a : _GEN_836; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_838 = 8'h46 == io_in_3 ? 8'h8c : _GEN_837; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_839 = 8'h47 == io_in_3 ? 8'h8e : _GEN_838; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_840 = 8'h48 == io_in_3 ? 8'h90 : _GEN_839; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_841 = 8'h49 == io_in_3 ? 8'h92 : _GEN_840; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_842 = 8'h4a == io_in_3 ? 8'h94 : _GEN_841; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_843 = 8'h4b == io_in_3 ? 8'h96 : _GEN_842; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_844 = 8'h4c == io_in_3 ? 8'h98 : _GEN_843; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_845 = 8'h4d == io_in_3 ? 8'h9a : _GEN_844; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_846 = 8'h4e == io_in_3 ? 8'h9c : _GEN_845; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_847 = 8'h4f == io_in_3 ? 8'h9e : _GEN_846; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_848 = 8'h50 == io_in_3 ? 8'ha0 : _GEN_847; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_849 = 8'h51 == io_in_3 ? 8'ha2 : _GEN_848; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_850 = 8'h52 == io_in_3 ? 8'ha4 : _GEN_849; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_851 = 8'h53 == io_in_3 ? 8'ha6 : _GEN_850; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_852 = 8'h54 == io_in_3 ? 8'ha8 : _GEN_851; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_853 = 8'h55 == io_in_3 ? 8'haa : _GEN_852; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_854 = 8'h56 == io_in_3 ? 8'hac : _GEN_853; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_855 = 8'h57 == io_in_3 ? 8'hae : _GEN_854; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_856 = 8'h58 == io_in_3 ? 8'hb0 : _GEN_855; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_857 = 8'h59 == io_in_3 ? 8'hb2 : _GEN_856; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_858 = 8'h5a == io_in_3 ? 8'hb4 : _GEN_857; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_859 = 8'h5b == io_in_3 ? 8'hb6 : _GEN_858; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_860 = 8'h5c == io_in_3 ? 8'hb8 : _GEN_859; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_861 = 8'h5d == io_in_3 ? 8'hba : _GEN_860; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_862 = 8'h5e == io_in_3 ? 8'hbc : _GEN_861; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_863 = 8'h5f == io_in_3 ? 8'hbe : _GEN_862; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_864 = 8'h60 == io_in_3 ? 8'hc0 : _GEN_863; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_865 = 8'h61 == io_in_3 ? 8'hc2 : _GEN_864; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_866 = 8'h62 == io_in_3 ? 8'hc4 : _GEN_865; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_867 = 8'h63 == io_in_3 ? 8'hc6 : _GEN_866; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_868 = 8'h64 == io_in_3 ? 8'hc8 : _GEN_867; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_869 = 8'h65 == io_in_3 ? 8'hca : _GEN_868; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_870 = 8'h66 == io_in_3 ? 8'hcc : _GEN_869; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_871 = 8'h67 == io_in_3 ? 8'hce : _GEN_870; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_872 = 8'h68 == io_in_3 ? 8'hd0 : _GEN_871; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_873 = 8'h69 == io_in_3 ? 8'hd2 : _GEN_872; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_874 = 8'h6a == io_in_3 ? 8'hd4 : _GEN_873; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_875 = 8'h6b == io_in_3 ? 8'hd6 : _GEN_874; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_876 = 8'h6c == io_in_3 ? 8'hd8 : _GEN_875; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_877 = 8'h6d == io_in_3 ? 8'hda : _GEN_876; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_878 = 8'h6e == io_in_3 ? 8'hdc : _GEN_877; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_879 = 8'h6f == io_in_3 ? 8'hde : _GEN_878; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_880 = 8'h70 == io_in_3 ? 8'he0 : _GEN_879; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_881 = 8'h71 == io_in_3 ? 8'he2 : _GEN_880; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_882 = 8'h72 == io_in_3 ? 8'he4 : _GEN_881; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_883 = 8'h73 == io_in_3 ? 8'he6 : _GEN_882; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_884 = 8'h74 == io_in_3 ? 8'he8 : _GEN_883; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_885 = 8'h75 == io_in_3 ? 8'hea : _GEN_884; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_886 = 8'h76 == io_in_3 ? 8'hec : _GEN_885; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_887 = 8'h77 == io_in_3 ? 8'hee : _GEN_886; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_888 = 8'h78 == io_in_3 ? 8'hf0 : _GEN_887; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_889 = 8'h79 == io_in_3 ? 8'hf2 : _GEN_888; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_890 = 8'h7a == io_in_3 ? 8'hf4 : _GEN_889; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_891 = 8'h7b == io_in_3 ? 8'hf6 : _GEN_890; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_892 = 8'h7c == io_in_3 ? 8'hf8 : _GEN_891; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_893 = 8'h7d == io_in_3 ? 8'hfa : _GEN_892; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_894 = 8'h7e == io_in_3 ? 8'hfc : _GEN_893; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_895 = 8'h7f == io_in_3 ? 8'hfe : _GEN_894; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_896 = 8'h80 == io_in_3 ? 8'h1b : _GEN_895; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_897 = 8'h81 == io_in_3 ? 8'h19 : _GEN_896; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_898 = 8'h82 == io_in_3 ? 8'h1f : _GEN_897; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_899 = 8'h83 == io_in_3 ? 8'h1d : _GEN_898; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_900 = 8'h84 == io_in_3 ? 8'h13 : _GEN_899; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_901 = 8'h85 == io_in_3 ? 8'h11 : _GEN_900; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_902 = 8'h86 == io_in_3 ? 8'h17 : _GEN_901; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_903 = 8'h87 == io_in_3 ? 8'h15 : _GEN_902; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_904 = 8'h88 == io_in_3 ? 8'hb : _GEN_903; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_905 = 8'h89 == io_in_3 ? 8'h9 : _GEN_904; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_906 = 8'h8a == io_in_3 ? 8'hf : _GEN_905; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_907 = 8'h8b == io_in_3 ? 8'hd : _GEN_906; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_908 = 8'h8c == io_in_3 ? 8'h3 : _GEN_907; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_909 = 8'h8d == io_in_3 ? 8'h1 : _GEN_908; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_910 = 8'h8e == io_in_3 ? 8'h7 : _GEN_909; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_911 = 8'h8f == io_in_3 ? 8'h5 : _GEN_910; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_912 = 8'h90 == io_in_3 ? 8'h3b : _GEN_911; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_913 = 8'h91 == io_in_3 ? 8'h39 : _GEN_912; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_914 = 8'h92 == io_in_3 ? 8'h3f : _GEN_913; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_915 = 8'h93 == io_in_3 ? 8'h3d : _GEN_914; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_916 = 8'h94 == io_in_3 ? 8'h33 : _GEN_915; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_917 = 8'h95 == io_in_3 ? 8'h31 : _GEN_916; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_918 = 8'h96 == io_in_3 ? 8'h37 : _GEN_917; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_919 = 8'h97 == io_in_3 ? 8'h35 : _GEN_918; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_920 = 8'h98 == io_in_3 ? 8'h2b : _GEN_919; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_921 = 8'h99 == io_in_3 ? 8'h29 : _GEN_920; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_922 = 8'h9a == io_in_3 ? 8'h2f : _GEN_921; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_923 = 8'h9b == io_in_3 ? 8'h2d : _GEN_922; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_924 = 8'h9c == io_in_3 ? 8'h23 : _GEN_923; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_925 = 8'h9d == io_in_3 ? 8'h21 : _GEN_924; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_926 = 8'h9e == io_in_3 ? 8'h27 : _GEN_925; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_927 = 8'h9f == io_in_3 ? 8'h25 : _GEN_926; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_928 = 8'ha0 == io_in_3 ? 8'h5b : _GEN_927; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_929 = 8'ha1 == io_in_3 ? 8'h59 : _GEN_928; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_930 = 8'ha2 == io_in_3 ? 8'h5f : _GEN_929; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_931 = 8'ha3 == io_in_3 ? 8'h5d : _GEN_930; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_932 = 8'ha4 == io_in_3 ? 8'h53 : _GEN_931; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_933 = 8'ha5 == io_in_3 ? 8'h51 : _GEN_932; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_934 = 8'ha6 == io_in_3 ? 8'h57 : _GEN_933; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_935 = 8'ha7 == io_in_3 ? 8'h55 : _GEN_934; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_936 = 8'ha8 == io_in_3 ? 8'h4b : _GEN_935; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_937 = 8'ha9 == io_in_3 ? 8'h49 : _GEN_936; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_938 = 8'haa == io_in_3 ? 8'h4f : _GEN_937; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_939 = 8'hab == io_in_3 ? 8'h4d : _GEN_938; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_940 = 8'hac == io_in_3 ? 8'h43 : _GEN_939; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_941 = 8'had == io_in_3 ? 8'h41 : _GEN_940; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_942 = 8'hae == io_in_3 ? 8'h47 : _GEN_941; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_943 = 8'haf == io_in_3 ? 8'h45 : _GEN_942; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_944 = 8'hb0 == io_in_3 ? 8'h7b : _GEN_943; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_945 = 8'hb1 == io_in_3 ? 8'h79 : _GEN_944; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_946 = 8'hb2 == io_in_3 ? 8'h7f : _GEN_945; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_947 = 8'hb3 == io_in_3 ? 8'h7d : _GEN_946; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_948 = 8'hb4 == io_in_3 ? 8'h73 : _GEN_947; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_949 = 8'hb5 == io_in_3 ? 8'h71 : _GEN_948; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_950 = 8'hb6 == io_in_3 ? 8'h77 : _GEN_949; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_951 = 8'hb7 == io_in_3 ? 8'h75 : _GEN_950; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_952 = 8'hb8 == io_in_3 ? 8'h6b : _GEN_951; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_953 = 8'hb9 == io_in_3 ? 8'h69 : _GEN_952; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_954 = 8'hba == io_in_3 ? 8'h6f : _GEN_953; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_955 = 8'hbb == io_in_3 ? 8'h6d : _GEN_954; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_956 = 8'hbc == io_in_3 ? 8'h63 : _GEN_955; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_957 = 8'hbd == io_in_3 ? 8'h61 : _GEN_956; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_958 = 8'hbe == io_in_3 ? 8'h67 : _GEN_957; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_959 = 8'hbf == io_in_3 ? 8'h65 : _GEN_958; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_960 = 8'hc0 == io_in_3 ? 8'h9b : _GEN_959; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_961 = 8'hc1 == io_in_3 ? 8'h99 : _GEN_960; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_962 = 8'hc2 == io_in_3 ? 8'h9f : _GEN_961; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_963 = 8'hc3 == io_in_3 ? 8'h9d : _GEN_962; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_964 = 8'hc4 == io_in_3 ? 8'h93 : _GEN_963; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_965 = 8'hc5 == io_in_3 ? 8'h91 : _GEN_964; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_966 = 8'hc6 == io_in_3 ? 8'h97 : _GEN_965; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_967 = 8'hc7 == io_in_3 ? 8'h95 : _GEN_966; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_968 = 8'hc8 == io_in_3 ? 8'h8b : _GEN_967; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_969 = 8'hc9 == io_in_3 ? 8'h89 : _GEN_968; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_970 = 8'hca == io_in_3 ? 8'h8f : _GEN_969; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_971 = 8'hcb == io_in_3 ? 8'h8d : _GEN_970; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_972 = 8'hcc == io_in_3 ? 8'h83 : _GEN_971; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_973 = 8'hcd == io_in_3 ? 8'h81 : _GEN_972; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_974 = 8'hce == io_in_3 ? 8'h87 : _GEN_973; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_975 = 8'hcf == io_in_3 ? 8'h85 : _GEN_974; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_976 = 8'hd0 == io_in_3 ? 8'hbb : _GEN_975; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_977 = 8'hd1 == io_in_3 ? 8'hb9 : _GEN_976; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_978 = 8'hd2 == io_in_3 ? 8'hbf : _GEN_977; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_979 = 8'hd3 == io_in_3 ? 8'hbd : _GEN_978; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_980 = 8'hd4 == io_in_3 ? 8'hb3 : _GEN_979; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_981 = 8'hd5 == io_in_3 ? 8'hb1 : _GEN_980; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_982 = 8'hd6 == io_in_3 ? 8'hb7 : _GEN_981; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_983 = 8'hd7 == io_in_3 ? 8'hb5 : _GEN_982; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_984 = 8'hd8 == io_in_3 ? 8'hab : _GEN_983; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_985 = 8'hd9 == io_in_3 ? 8'ha9 : _GEN_984; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_986 = 8'hda == io_in_3 ? 8'haf : _GEN_985; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_987 = 8'hdb == io_in_3 ? 8'had : _GEN_986; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_988 = 8'hdc == io_in_3 ? 8'ha3 : _GEN_987; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_989 = 8'hdd == io_in_3 ? 8'ha1 : _GEN_988; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_990 = 8'hde == io_in_3 ? 8'ha7 : _GEN_989; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_991 = 8'hdf == io_in_3 ? 8'ha5 : _GEN_990; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_992 = 8'he0 == io_in_3 ? 8'hdb : _GEN_991; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_993 = 8'he1 == io_in_3 ? 8'hd9 : _GEN_992; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_994 = 8'he2 == io_in_3 ? 8'hdf : _GEN_993; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_995 = 8'he3 == io_in_3 ? 8'hdd : _GEN_994; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_996 = 8'he4 == io_in_3 ? 8'hd3 : _GEN_995; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_997 = 8'he5 == io_in_3 ? 8'hd1 : _GEN_996; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_998 = 8'he6 == io_in_3 ? 8'hd7 : _GEN_997; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_999 = 8'he7 == io_in_3 ? 8'hd5 : _GEN_998; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1000 = 8'he8 == io_in_3 ? 8'hcb : _GEN_999; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1001 = 8'he9 == io_in_3 ? 8'hc9 : _GEN_1000; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1002 = 8'hea == io_in_3 ? 8'hcf : _GEN_1001; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1003 = 8'heb == io_in_3 ? 8'hcd : _GEN_1002; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1004 = 8'hec == io_in_3 ? 8'hc3 : _GEN_1003; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1005 = 8'hed == io_in_3 ? 8'hc1 : _GEN_1004; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1006 = 8'hee == io_in_3 ? 8'hc7 : _GEN_1005; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1007 = 8'hef == io_in_3 ? 8'hc5 : _GEN_1006; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1008 = 8'hf0 == io_in_3 ? 8'hfb : _GEN_1007; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1009 = 8'hf1 == io_in_3 ? 8'hf9 : _GEN_1008; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1010 = 8'hf2 == io_in_3 ? 8'hff : _GEN_1009; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1011 = 8'hf3 == io_in_3 ? 8'hfd : _GEN_1010; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1012 = 8'hf4 == io_in_3 ? 8'hf3 : _GEN_1011; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1013 = 8'hf5 == io_in_3 ? 8'hf1 : _GEN_1012; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1014 = 8'hf6 == io_in_3 ? 8'hf7 : _GEN_1013; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1015 = 8'hf7 == io_in_3 ? 8'hf5 : _GEN_1014; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1016 = 8'hf8 == io_in_3 ? 8'heb : _GEN_1015; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1017 = 8'hf9 == io_in_3 ? 8'he9 : _GEN_1016; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1018 = 8'hfa == io_in_3 ? 8'hef : _GEN_1017; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1019 = 8'hfb == io_in_3 ? 8'hed : _GEN_1018; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1020 = 8'hfc == io_in_3 ? 8'he3 : _GEN_1019; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1021 = 8'hfd == io_in_3 ? 8'he1 : _GEN_1020; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1022 = 8'hfe == io_in_3 ? 8'he7 : _GEN_1021; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _GEN_1023 = 8'hff == io_in_3 ? 8'he5 : _GEN_1022; // @[AES_PipelinedElasticBuffer.scala 330:53 AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _T_10 = _T_9 ^ _GEN_1023; // @[AES_PipelinedElasticBuffer.scala 330:53]
  wire [7:0] _T_12 = _GEN_255 ^ io_in_0; // @[AES_PipelinedElasticBuffer.scala 331:31]
  wire [7:0] _T_13 = _T_12 ^ io_in_1; // @[AES_PipelinedElasticBuffer.scala 331:42]
  wire [7:0] _T_14 = _T_13 ^ io_in_2; // @[AES_PipelinedElasticBuffer.scala 331:53]
  assign io_out_0 = _T_2 ^ io_in_3; // @[AES_PipelinedElasticBuffer.scala 328:70]
  assign io_out_1 = _T_6 ^ io_in_3; // @[AES_PipelinedElasticBuffer.scala 329:70]
  assign io_out_2 = _T_10 ^ io_in_3; // @[AES_PipelinedElasticBuffer.scala 330:70]
  assign io_out_3 = _T_14 ^ _GEN_1023; // @[AES_PipelinedElasticBuffer.scala 331:64]
endmodule
module AES_MixColumns(
  output [7:0] io_out_state_0_0,
  output [7:0] io_out_state_0_1,
  output [7:0] io_out_state_0_2,
  output [7:0] io_out_state_0_3,
  output [7:0] io_out_state_1_0,
  output [7:0] io_out_state_1_1,
  output [7:0] io_out_state_1_2,
  output [7:0] io_out_state_1_3,
  output [7:0] io_out_state_2_0,
  output [7:0] io_out_state_2_1,
  output [7:0] io_out_state_2_2,
  output [7:0] io_out_state_2_3,
  output [7:0] io_out_state_3_0,
  output [7:0] io_out_state_3_1,
  output [7:0] io_out_state_3_2,
  output [7:0] io_out_state_3_3,
  input  [7:0] io_in_state_0_0,
  input  [7:0] io_in_state_0_1,
  input  [7:0] io_in_state_0_2,
  input  [7:0] io_in_state_0_3,
  input  [7:0] io_in_state_1_0,
  input  [7:0] io_in_state_1_1,
  input  [7:0] io_in_state_1_2,
  input  [7:0] io_in_state_1_3,
  input  [7:0] io_in_state_2_0,
  input  [7:0] io_in_state_2_1,
  input  [7:0] io_in_state_2_2,
  input  [7:0] io_in_state_2_3,
  input  [7:0] io_in_state_3_0,
  input  [7:0] io_in_state_3_1,
  input  [7:0] io_in_state_3_2,
  input  [7:0] io_in_state_3_3
);
  wire [7:0] PEs_0_io_in_0; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_0_io_in_1; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_0_io_in_2; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_0_io_in_3; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_0_io_out_0; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_0_io_out_1; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_0_io_out_2; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_0_io_out_3; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_1_io_in_0; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_1_io_in_1; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_1_io_in_2; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_1_io_in_3; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_1_io_out_0; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_1_io_out_1; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_1_io_out_2; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_1_io_out_3; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_2_io_in_0; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_2_io_in_1; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_2_io_in_2; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_2_io_in_3; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_2_io_out_0; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_2_io_out_1; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_2_io_out_2; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_2_io_out_3; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_3_io_in_0; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_3_io_in_1; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_3_io_in_2; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_3_io_in_3; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_3_io_out_0; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_3_io_out_1; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_3_io_out_2; // @[AES_PipelinedElasticBuffer.scala 278:20]
  wire [7:0] PEs_3_io_out_3; // @[AES_PipelinedElasticBuffer.scala 278:20]
  AES_MixColumn PEs_0 ( // @[AES_PipelinedElasticBuffer.scala 278:20]
    .io_in_0(PEs_0_io_in_0),
    .io_in_1(PEs_0_io_in_1),
    .io_in_2(PEs_0_io_in_2),
    .io_in_3(PEs_0_io_in_3),
    .io_out_0(PEs_0_io_out_0),
    .io_out_1(PEs_0_io_out_1),
    .io_out_2(PEs_0_io_out_2),
    .io_out_3(PEs_0_io_out_3)
  );
  AES_MixColumn PEs_1 ( // @[AES_PipelinedElasticBuffer.scala 278:20]
    .io_in_0(PEs_1_io_in_0),
    .io_in_1(PEs_1_io_in_1),
    .io_in_2(PEs_1_io_in_2),
    .io_in_3(PEs_1_io_in_3),
    .io_out_0(PEs_1_io_out_0),
    .io_out_1(PEs_1_io_out_1),
    .io_out_2(PEs_1_io_out_2),
    .io_out_3(PEs_1_io_out_3)
  );
  AES_MixColumn PEs_2 ( // @[AES_PipelinedElasticBuffer.scala 278:20]
    .io_in_0(PEs_2_io_in_0),
    .io_in_1(PEs_2_io_in_1),
    .io_in_2(PEs_2_io_in_2),
    .io_in_3(PEs_2_io_in_3),
    .io_out_0(PEs_2_io_out_0),
    .io_out_1(PEs_2_io_out_1),
    .io_out_2(PEs_2_io_out_2),
    .io_out_3(PEs_2_io_out_3)
  );
  AES_MixColumn PEs_3 ( // @[AES_PipelinedElasticBuffer.scala 278:20]
    .io_in_0(PEs_3_io_in_0),
    .io_in_1(PEs_3_io_in_1),
    .io_in_2(PEs_3_io_in_2),
    .io_in_3(PEs_3_io_in_3),
    .io_out_0(PEs_3_io_out_0),
    .io_out_1(PEs_3_io_out_1),
    .io_out_2(PEs_3_io_out_2),
    .io_out_3(PEs_3_io_out_3)
  );
  assign io_out_state_0_0 = PEs_0_io_out_0; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_0_1 = PEs_0_io_out_1; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_0_2 = PEs_0_io_out_2; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_0_3 = PEs_0_io_out_3; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_1_0 = PEs_1_io_out_0; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_1_1 = PEs_1_io_out_1; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_1_2 = PEs_1_io_out_2; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_1_3 = PEs_1_io_out_3; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_2_0 = PEs_2_io_out_0; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_2_1 = PEs_2_io_out_1; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_2_2 = PEs_2_io_out_2; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_2_3 = PEs_2_io_out_3; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_3_0 = PEs_3_io_out_0; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_3_1 = PEs_3_io_out_1; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_3_2 = PEs_3_io_out_2; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign io_out_state_3_3 = PEs_3_io_out_3; // @[AES_PipelinedElasticBuffer.scala 285:21]
  assign PEs_0_io_in_0 = io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_0_io_in_1 = io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_0_io_in_2 = io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_0_io_in_3 = io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_1_io_in_0 = io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_1_io_in_1 = io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_1_io_in_2 = io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_1_io_in_3 = io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_2_io_in_0 = io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_2_io_in_1 = io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_2_io_in_2 = io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_2_io_in_3 = io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_3_io_in_0 = io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_3_io_in_1 = io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_3_io_in_2 = io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 284:18]
  assign PEs_3_io_in_3 = io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 284:18]
endmodule
module AES_RotWord(
  output [31:0] io_out,
  input  [31:0] io_in
);
  wire [23:0] hi = io_in[23:0]; // @[AES_PipelinedElasticBuffer.scala 266:22]
  wire [7:0] lo = io_in[31:24]; // @[AES_PipelinedElasticBuffer.scala 266:35]
  assign io_out = {hi,lo}; // @[Cat.scala 30:58]
endmodule
module AES_SubWord(
  output [31:0] io_out,
  input  [31:0] io_in
);
  wire [7:0] PEs_0_io_in; // @[AES_PipelinedElasticBuffer.scala 252:20]
  wire [7:0] PEs_0_io_out; // @[AES_PipelinedElasticBuffer.scala 252:20]
  wire [7:0] PEs_1_io_in; // @[AES_PipelinedElasticBuffer.scala 252:20]
  wire [7:0] PEs_1_io_out; // @[AES_PipelinedElasticBuffer.scala 252:20]
  wire [7:0] PEs_2_io_in; // @[AES_PipelinedElasticBuffer.scala 252:20]
  wire [7:0] PEs_2_io_out; // @[AES_PipelinedElasticBuffer.scala 252:20]
  wire [7:0] PEs_3_io_in; // @[AES_PipelinedElasticBuffer.scala 252:20]
  wire [7:0] PEs_3_io_out; // @[AES_PipelinedElasticBuffer.scala 252:20]
  wire [15:0] lo = {PEs_1_io_out,PEs_0_io_out}; // @[Cat.scala 30:58]
  wire [15:0] hi = {PEs_3_io_out,PEs_2_io_out}; // @[Cat.scala 30:58]
  AES_S PEs_0 ( // @[AES_PipelinedElasticBuffer.scala 252:20]
    .io_in(PEs_0_io_in),
    .io_out(PEs_0_io_out)
  );
  AES_S PEs_1 ( // @[AES_PipelinedElasticBuffer.scala 252:20]
    .io_in(PEs_1_io_in),
    .io_out(PEs_1_io_out)
  );
  AES_S PEs_2 ( // @[AES_PipelinedElasticBuffer.scala 252:20]
    .io_in(PEs_2_io_in),
    .io_out(PEs_2_io_out)
  );
  AES_S PEs_3 ( // @[AES_PipelinedElasticBuffer.scala 252:20]
    .io_in(PEs_3_io_in),
    .io_out(PEs_3_io_out)
  );
  assign io_out = {hi,lo}; // @[Cat.scala 30:58]
  assign PEs_0_io_in = io_in[7:0]; // @[AES_PipelinedElasticBuffer.scala 253:22]
  assign PEs_1_io_in = io_in[15:8]; // @[AES_PipelinedElasticBuffer.scala 253:22]
  assign PEs_2_io_in = io_in[23:16]; // @[AES_PipelinedElasticBuffer.scala 253:22]
  assign PEs_3_io_in = io_in[31:24]; // @[AES_PipelinedElasticBuffer.scala 253:22]
endmodule
module AES_GetNewKey(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_4 = sub_io_out ^ 32'h1000000; // @[AES_PipelinedElasticBuffer.scala 232:20]
  wire [31:0] w5 = _T_4 ^ w0; // @[AES_PipelinedElasticBuffer.scala 232:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_PipelinedElasticBuffer.scala 233:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_PipelinedElasticBuffer.scala 234:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_PipelinedElasticBuffer.scala 235:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 211:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 214:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 215:13]
endmodule
module AES_ProcessingElement(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 149:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 150:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 150:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:23 AES_PipelinedElasticBuffer.scala 158:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 165:21 AES_PipelinedElasticBuffer.scala 165:21]
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 171:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_PipelinedElasticBuffer.scala 179:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_PipelinedElasticBuffer.scala 182:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey key ( // @[AES_PipelinedElasticBuffer.scala 191:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 153:27]
  assign io_out_bits_state_0_0 = mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_1 = mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_2 = mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_3 = mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_0 = mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_1 = mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_2 = mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_3 = mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_0 = mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_1 = mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_2 = mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_3 = mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_0 = mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_1 = mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_2 = mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_3 = mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_0 = key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_1 = key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_2 = key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_3 = key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_0 = key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_1 = key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_2 = key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_3 = key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_0 = key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_1 = key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_2 = key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_3 = key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_0 = key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_1 = key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_2 = key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_3 = key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 152:18]
  assign sub_io_in_state_0_0 = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_1 = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_2 = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_3 = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_0 = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_1 = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_2 = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_3 = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_0 = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_1 = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_2 = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_3 = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_0 = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_1 = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_2 = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_3 = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign key_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 167:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 149:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 149:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 161:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_1(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_4 = sub_io_out ^ 32'h2000000; // @[AES_PipelinedElasticBuffer.scala 232:20]
  wire [31:0] w5 = _T_4 ^ w0; // @[AES_PipelinedElasticBuffer.scala 232:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_PipelinedElasticBuffer.scala 233:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_PipelinedElasticBuffer.scala 234:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_PipelinedElasticBuffer.scala 235:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 211:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 214:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 215:13]
endmodule
module AES_ProcessingElement_1(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 149:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 150:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 150:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:23 AES_PipelinedElasticBuffer.scala 158:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 165:21 AES_PipelinedElasticBuffer.scala 165:21]
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 171:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_PipelinedElasticBuffer.scala 179:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_PipelinedElasticBuffer.scala 182:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey_1 key ( // @[AES_PipelinedElasticBuffer.scala 191:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 153:27]
  assign io_out_bits_state_0_0 = mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_1 = mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_2 = mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_3 = mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_0 = mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_1 = mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_2 = mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_3 = mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_0 = mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_1 = mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_2 = mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_3 = mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_0 = mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_1 = mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_2 = mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_3 = mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_0 = key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_1 = key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_2 = key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_3 = key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_0 = key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_1 = key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_2 = key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_3 = key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_0 = key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_1 = key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_2 = key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_3 = key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_0 = key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_1 = key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_2 = key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_3 = key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 152:18]
  assign sub_io_in_state_0_0 = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_1 = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_2 = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_3 = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_0 = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_1 = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_2 = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_3 = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_0 = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_1 = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_2 = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_3 = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_0 = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_1 = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_2 = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_3 = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign key_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 167:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 149:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 149:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 161:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_2(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_4 = sub_io_out ^ 32'h4000000; // @[AES_PipelinedElasticBuffer.scala 232:20]
  wire [31:0] w5 = _T_4 ^ w0; // @[AES_PipelinedElasticBuffer.scala 232:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_PipelinedElasticBuffer.scala 233:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_PipelinedElasticBuffer.scala 234:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_PipelinedElasticBuffer.scala 235:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 211:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 214:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 215:13]
endmodule
module AES_ProcessingElement_2(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 149:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 150:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 150:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:23 AES_PipelinedElasticBuffer.scala 158:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 165:21 AES_PipelinedElasticBuffer.scala 165:21]
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 171:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_PipelinedElasticBuffer.scala 179:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_PipelinedElasticBuffer.scala 182:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey_2 key ( // @[AES_PipelinedElasticBuffer.scala 191:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 153:27]
  assign io_out_bits_state_0_0 = mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_1 = mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_2 = mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_3 = mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_0 = mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_1 = mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_2 = mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_3 = mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_0 = mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_1 = mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_2 = mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_3 = mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_0 = mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_1 = mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_2 = mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_3 = mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_0 = key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_1 = key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_2 = key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_3 = key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_0 = key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_1 = key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_2 = key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_3 = key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_0 = key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_1 = key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_2 = key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_3 = key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_0 = key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_1 = key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_2 = key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_3 = key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 152:18]
  assign sub_io_in_state_0_0 = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_1 = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_2 = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_3 = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_0 = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_1 = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_2 = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_3 = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_0 = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_1 = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_2 = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_3 = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_0 = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_1 = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_2 = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_3 = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign key_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 167:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 149:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 149:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 161:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_3(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_4 = sub_io_out ^ 32'h8000000; // @[AES_PipelinedElasticBuffer.scala 232:20]
  wire [31:0] w5 = _T_4 ^ w0; // @[AES_PipelinedElasticBuffer.scala 232:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_PipelinedElasticBuffer.scala 233:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_PipelinedElasticBuffer.scala 234:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_PipelinedElasticBuffer.scala 235:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 211:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 214:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 215:13]
endmodule
module AES_ProcessingElement_3(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 149:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 150:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 150:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:23 AES_PipelinedElasticBuffer.scala 158:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 165:21 AES_PipelinedElasticBuffer.scala 165:21]
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 171:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_PipelinedElasticBuffer.scala 179:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_PipelinedElasticBuffer.scala 182:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey_3 key ( // @[AES_PipelinedElasticBuffer.scala 191:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 153:27]
  assign io_out_bits_state_0_0 = mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_1 = mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_2 = mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_3 = mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_0 = mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_1 = mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_2 = mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_3 = mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_0 = mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_1 = mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_2 = mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_3 = mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_0 = mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_1 = mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_2 = mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_3 = mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_0 = key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_1 = key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_2 = key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_3 = key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_0 = key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_1 = key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_2 = key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_3 = key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_0 = key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_1 = key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_2 = key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_3 = key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_0 = key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_1 = key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_2 = key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_3 = key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 152:18]
  assign sub_io_in_state_0_0 = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_1 = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_2 = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_3 = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_0 = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_1 = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_2 = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_3 = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_0 = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_1 = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_2 = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_3 = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_0 = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_1 = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_2 = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_3 = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign key_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 167:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 149:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 149:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 161:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_4(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_4 = sub_io_out ^ 32'h10000000; // @[AES_PipelinedElasticBuffer.scala 232:20]
  wire [31:0] w5 = _T_4 ^ w0; // @[AES_PipelinedElasticBuffer.scala 232:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_PipelinedElasticBuffer.scala 233:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_PipelinedElasticBuffer.scala 234:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_PipelinedElasticBuffer.scala 235:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 211:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 214:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 215:13]
endmodule
module AES_ProcessingElement_4(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 149:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 150:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 150:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:23 AES_PipelinedElasticBuffer.scala 158:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 165:21 AES_PipelinedElasticBuffer.scala 165:21]
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 171:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_PipelinedElasticBuffer.scala 179:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_PipelinedElasticBuffer.scala 182:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey_4 key ( // @[AES_PipelinedElasticBuffer.scala 191:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 153:27]
  assign io_out_bits_state_0_0 = mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_1 = mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_2 = mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_3 = mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_0 = mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_1 = mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_2 = mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_3 = mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_0 = mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_1 = mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_2 = mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_3 = mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_0 = mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_1 = mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_2 = mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_3 = mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_0 = key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_1 = key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_2 = key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_3 = key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_0 = key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_1 = key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_2 = key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_3 = key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_0 = key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_1 = key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_2 = key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_3 = key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_0 = key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_1 = key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_2 = key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_3 = key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 152:18]
  assign sub_io_in_state_0_0 = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_1 = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_2 = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_3 = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_0 = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_1 = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_2 = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_3 = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_0 = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_1 = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_2 = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_3 = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_0 = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_1 = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_2 = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_3 = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign key_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 167:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 149:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 149:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 161:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_5(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_4 = sub_io_out ^ 32'h20000000; // @[AES_PipelinedElasticBuffer.scala 232:20]
  wire [31:0] w5 = _T_4 ^ w0; // @[AES_PipelinedElasticBuffer.scala 232:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_PipelinedElasticBuffer.scala 233:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_PipelinedElasticBuffer.scala 234:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_PipelinedElasticBuffer.scala 235:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 211:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 214:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 215:13]
endmodule
module AES_ProcessingElement_5(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 149:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 150:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 150:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:23 AES_PipelinedElasticBuffer.scala 158:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 165:21 AES_PipelinedElasticBuffer.scala 165:21]
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 171:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_PipelinedElasticBuffer.scala 179:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_PipelinedElasticBuffer.scala 182:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey_5 key ( // @[AES_PipelinedElasticBuffer.scala 191:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 153:27]
  assign io_out_bits_state_0_0 = mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_1 = mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_2 = mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_3 = mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_0 = mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_1 = mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_2 = mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_3 = mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_0 = mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_1 = mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_2 = mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_3 = mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_0 = mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_1 = mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_2 = mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_3 = mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_0 = key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_1 = key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_2 = key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_3 = key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_0 = key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_1 = key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_2 = key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_3 = key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_0 = key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_1 = key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_2 = key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_3 = key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_0 = key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_1 = key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_2 = key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_3 = key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 152:18]
  assign sub_io_in_state_0_0 = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_1 = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_2 = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_3 = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_0 = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_1 = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_2 = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_3 = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_0 = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_1 = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_2 = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_3 = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_0 = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_1 = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_2 = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_3 = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign key_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 167:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 149:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 149:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 161:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_6(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_4 = sub_io_out ^ 32'h40000000; // @[AES_PipelinedElasticBuffer.scala 232:20]
  wire [31:0] w5 = _T_4 ^ w0; // @[AES_PipelinedElasticBuffer.scala 232:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_PipelinedElasticBuffer.scala 233:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_PipelinedElasticBuffer.scala 234:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_PipelinedElasticBuffer.scala 235:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 211:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 214:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 215:13]
endmodule
module AES_ProcessingElement_6(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 149:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 150:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 150:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:23 AES_PipelinedElasticBuffer.scala 158:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 165:21 AES_PipelinedElasticBuffer.scala 165:21]
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 171:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_PipelinedElasticBuffer.scala 179:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_PipelinedElasticBuffer.scala 182:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey_6 key ( // @[AES_PipelinedElasticBuffer.scala 191:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 153:27]
  assign io_out_bits_state_0_0 = mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_1 = mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_2 = mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_3 = mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_0 = mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_1 = mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_2 = mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_3 = mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_0 = mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_1 = mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_2 = mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_3 = mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_0 = mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_1 = mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_2 = mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_3 = mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_0 = key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_1 = key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_2 = key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_3 = key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_0 = key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_1 = key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_2 = key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_3 = key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_0 = key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_1 = key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_2 = key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_3 = key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_0 = key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_1 = key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_2 = key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_3 = key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 152:18]
  assign sub_io_in_state_0_0 = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_1 = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_2 = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_3 = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_0 = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_1 = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_2 = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_3 = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_0 = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_1 = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_2 = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_3 = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_0 = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_1 = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_2 = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_3 = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign key_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 167:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 149:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 149:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 161:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_7(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_4 = sub_io_out ^ 32'h80000000; // @[AES_PipelinedElasticBuffer.scala 232:20]
  wire [31:0] w5 = _T_4 ^ w0; // @[AES_PipelinedElasticBuffer.scala 232:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_PipelinedElasticBuffer.scala 233:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_PipelinedElasticBuffer.scala 234:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_PipelinedElasticBuffer.scala 235:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 211:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 214:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 215:13]
endmodule
module AES_ProcessingElement_7(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 149:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 150:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 150:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:23 AES_PipelinedElasticBuffer.scala 158:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 165:21 AES_PipelinedElasticBuffer.scala 165:21]
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 171:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_PipelinedElasticBuffer.scala 179:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_PipelinedElasticBuffer.scala 182:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey_7 key ( // @[AES_PipelinedElasticBuffer.scala 191:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 153:27]
  assign io_out_bits_state_0_0 = mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_1 = mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_2 = mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_3 = mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_0 = mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_1 = mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_2 = mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_3 = mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_0 = mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_1 = mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_2 = mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_3 = mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_0 = mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_1 = mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_2 = mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_3 = mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_0 = key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_1 = key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_2 = key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_3 = key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_0 = key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_1 = key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_2 = key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_3 = key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_0 = key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_1 = key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_2 = key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_3 = key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_0 = key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_1 = key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_2 = key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_3 = key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 152:18]
  assign sub_io_in_state_0_0 = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_1 = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_2 = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_3 = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_0 = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_1 = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_2 = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_3 = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_0 = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_1 = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_2 = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_3 = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_0 = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_1 = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_2 = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_3 = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign key_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 167:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 149:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 149:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 161:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_8(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_4 = sub_io_out ^ 32'h1b000000; // @[AES_PipelinedElasticBuffer.scala 232:20]
  wire [31:0] w5 = _T_4 ^ w0; // @[AES_PipelinedElasticBuffer.scala 232:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_PipelinedElasticBuffer.scala 233:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_PipelinedElasticBuffer.scala 234:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_PipelinedElasticBuffer.scala 235:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 211:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 214:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 215:13]
endmodule
module AES_ProcessingElement_8(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 149:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 150:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 150:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:23 AES_PipelinedElasticBuffer.scala 158:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 165:21 AES_PipelinedElasticBuffer.scala 165:21]
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 171:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_PipelinedElasticBuffer.scala 179:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_PipelinedElasticBuffer.scala 182:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey_8 key ( // @[AES_PipelinedElasticBuffer.scala 191:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 153:27]
  assign io_out_bits_state_0_0 = mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_1 = mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_2 = mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_3 = mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_0 = mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_1 = mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_2 = mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_3 = mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_0 = mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_1 = mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_2 = mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_3 = mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_0 = mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_1 = mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_2 = mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_3 = mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_0 = key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_1 = key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_2 = key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_3 = key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_0 = key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_1 = key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_2 = key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_3 = key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_0 = key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_1 = key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_2 = key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_3 = key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_0 = key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_1 = key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_2 = key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_3 = key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 152:18]
  assign sub_io_in_state_0_0 = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_1 = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_2 = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_3 = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_0 = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_1 = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_2 = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_3 = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_0 = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_1 = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_2 = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_3 = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_0 = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_1 = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_2 = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_3 = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign key_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 167:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 149:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 149:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 161:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_GetNewKey_9(
  output [7:0] io_out_key_0_0,
  output [7:0] io_out_key_0_1,
  output [7:0] io_out_key_0_2,
  output [7:0] io_out_key_0_3,
  output [7:0] io_out_key_1_0,
  output [7:0] io_out_key_1_1,
  output [7:0] io_out_key_1_2,
  output [7:0] io_out_key_1_3,
  output [7:0] io_out_key_2_0,
  output [7:0] io_out_key_2_1,
  output [7:0] io_out_key_2_2,
  output [7:0] io_out_key_2_3,
  output [7:0] io_out_key_3_0,
  output [7:0] io_out_key_3_1,
  output [7:0] io_out_key_3_2,
  output [7:0] io_out_key_3_3,
  input  [7:0] io_in_key_0_0,
  input  [7:0] io_in_key_0_1,
  input  [7:0] io_in_key_0_2,
  input  [7:0] io_in_key_0_3,
  input  [7:0] io_in_key_1_0,
  input  [7:0] io_in_key_1_1,
  input  [7:0] io_in_key_1_2,
  input  [7:0] io_in_key_1_3,
  input  [7:0] io_in_key_2_0,
  input  [7:0] io_in_key_2_1,
  input  [7:0] io_in_key_2_2,
  input  [7:0] io_in_key_2_3,
  input  [7:0] io_in_key_3_0,
  input  [7:0] io_in_key_3_1,
  input  [7:0] io_in_key_3_2,
  input  [7:0] io_in_key_3_3
);
  wire [31:0] rot_io_out; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] rot_io_in; // @[AES_PipelinedElasticBuffer.scala 211:19]
  wire [31:0] sub_io_out; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] sub_io_in; // @[AES_PipelinedElasticBuffer.scala 214:19]
  wire [31:0] w0 = {io_in_key_0_0,io_in_key_0_1,io_in_key_0_2,io_in_key_0_3}; // @[Cat.scala 30:58]
  wire [31:0] w1 = {io_in_key_1_0,io_in_key_1_1,io_in_key_1_2,io_in_key_1_3}; // @[Cat.scala 30:58]
  wire [31:0] w2 = {io_in_key_2_0,io_in_key_2_1,io_in_key_2_2,io_in_key_2_3}; // @[Cat.scala 30:58]
  wire [15:0] lo_3 = {io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = {io_in_key_3_0,io_in_key_3_1}; // @[Cat.scala 30:58]
  wire [31:0] w3 = {io_in_key_3_0,io_in_key_3_1,io_in_key_3_2,io_in_key_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_4 = sub_io_out ^ 32'h36000000; // @[AES_PipelinedElasticBuffer.scala 232:20]
  wire [31:0] w5 = _T_4 ^ w0; // @[AES_PipelinedElasticBuffer.scala 232:27]
  wire [31:0] w6 = w5 ^ w1; // @[AES_PipelinedElasticBuffer.scala 233:12]
  wire [31:0] w7 = w6 ^ w2; // @[AES_PipelinedElasticBuffer.scala 234:12]
  wire [31:0] w8 = w7 ^ w3; // @[AES_PipelinedElasticBuffer.scala 235:12]
  AES_RotWord rot ( // @[AES_PipelinedElasticBuffer.scala 211:19]
    .io_out(rot_io_out),
    .io_in(rot_io_in)
  );
  AES_SubWord sub ( // @[AES_PipelinedElasticBuffer.scala 214:19]
    .io_out(sub_io_out),
    .io_in(sub_io_in)
  );
  assign io_out_key_0_0 = w5[31:24]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_1 = w5[23:16]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_2 = w5[15:8]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_0_3 = w5[7:0]; // @[AES_PipelinedElasticBuffer.scala 238:29]
  assign io_out_key_1_0 = w6[31:24]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_1 = w6[23:16]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_2 = w6[15:8]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_1_3 = w6[7:0]; // @[AES_PipelinedElasticBuffer.scala 239:29]
  assign io_out_key_2_0 = w7[31:24]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_1 = w7[23:16]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_2 = w7[15:8]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_2_3 = w7[7:0]; // @[AES_PipelinedElasticBuffer.scala 240:29]
  assign io_out_key_3_0 = w8[31:24]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_1 = w8[23:16]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_2 = w8[15:8]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign io_out_key_3_3 = w8[7:0]; // @[AES_PipelinedElasticBuffer.scala 241:29]
  assign rot_io_in = {hi_3,lo_3}; // @[Cat.scala 30:58]
  assign sub_io_in = rot_io_out; // @[AES_PipelinedElasticBuffer.scala 215:13]
endmodule
module AES_ProcessingElement_9(
  input        clock,
  input        reset,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits_state_0_0,
  output [7:0] io_out_bits_state_0_1,
  output [7:0] io_out_bits_state_0_2,
  output [7:0] io_out_bits_state_0_3,
  output [7:0] io_out_bits_state_1_0,
  output [7:0] io_out_bits_state_1_1,
  output [7:0] io_out_bits_state_1_2,
  output [7:0] io_out_bits_state_1_3,
  output [7:0] io_out_bits_state_2_0,
  output [7:0] io_out_bits_state_2_1,
  output [7:0] io_out_bits_state_2_2,
  output [7:0] io_out_bits_state_2_3,
  output [7:0] io_out_bits_state_3_0,
  output [7:0] io_out_bits_state_3_1,
  output [7:0] io_out_bits_state_3_2,
  output [7:0] io_out_bits_state_3_3,
  output [7:0] io_out_bits_key_0_0,
  output [7:0] io_out_bits_key_0_1,
  output [7:0] io_out_bits_key_0_2,
  output [7:0] io_out_bits_key_0_3,
  output [7:0] io_out_bits_key_1_0,
  output [7:0] io_out_bits_key_1_1,
  output [7:0] io_out_bits_key_1_2,
  output [7:0] io_out_bits_key_1_3,
  output [7:0] io_out_bits_key_2_0,
  output [7:0] io_out_bits_key_2_1,
  output [7:0] io_out_bits_key_2_2,
  output [7:0] io_out_bits_key_2_3,
  output [7:0] io_out_bits_key_3_0,
  output [7:0] io_out_bits_key_3_1,
  output [7:0] io_out_bits_key_3_2,
  output [7:0] io_out_bits_key_3_3,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits_state_0_0,
  input  [7:0] io_in_bits_state_0_1,
  input  [7:0] io_in_bits_state_0_2,
  input  [7:0] io_in_bits_state_0_3,
  input  [7:0] io_in_bits_state_1_0,
  input  [7:0] io_in_bits_state_1_1,
  input  [7:0] io_in_bits_state_1_2,
  input  [7:0] io_in_bits_state_1_3,
  input  [7:0] io_in_bits_state_2_0,
  input  [7:0] io_in_bits_state_2_1,
  input  [7:0] io_in_bits_state_2_2,
  input  [7:0] io_in_bits_state_2_3,
  input  [7:0] io_in_bits_state_3_0,
  input  [7:0] io_in_bits_state_3_1,
  input  [7:0] io_in_bits_state_3_2,
  input  [7:0] io_in_bits_state_3_3,
  input  [7:0] io_in_bits_key_0_0,
  input  [7:0] io_in_bits_key_0_1,
  input  [7:0] io_in_bits_key_0_2,
  input  [7:0] io_in_bits_key_0_3,
  input  [7:0] io_in_bits_key_1_0,
  input  [7:0] io_in_bits_key_1_1,
  input  [7:0] io_in_bits_key_1_2,
  input  [7:0] io_in_bits_key_1_3,
  input  [7:0] io_in_bits_key_2_0,
  input  [7:0] io_in_bits_key_2_1,
  input  [7:0] io_in_bits_key_2_2,
  input  [7:0] io_in_bits_key_2_3,
  input  [7:0] io_in_bits_key_3_0,
  input  [7:0] io_in_bits_key_3_1,
  input  [7:0] io_in_bits_key_3_2,
  input  [7:0] io_in_bits_key_3_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] sub_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 171:19]
  wire [7:0] shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] shift_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 179:21]
  wire [7:0] mix_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_0_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_1_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_2_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_0; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_1; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_2; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] mix_io_in_state_3_3; // @[AES_PipelinedElasticBuffer.scala 182:19]
  wire [7:0] key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_0_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_1_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_2_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_0; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_1; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_2; // @[AES_PipelinedElasticBuffer.scala 191:19]
  wire [7:0] key_io_in_key_3_3; // @[AES_PipelinedElasticBuffer.scala 191:19]
  reg [7:0] data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_state_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_0_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_1_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_2_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_0; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_1; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_2; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg [7:0] data_1_key_3_3; // @[AES_PipelinedElasticBuffer.scala 147:21]
  reg  head; // @[AES_PipelinedElasticBuffer.scala 148:21]
  reg  tail; // @[AES_PipelinedElasticBuffer.scala 149:21]
  reg  full_0; // @[AES_PipelinedElasticBuffer.scala 150:21]
  reg  full_1; // @[AES_PipelinedElasticBuffer.scala 150:21]
  wire [7:0] input_state_0_0 = head ? data_1_state_0_0 : data_0_state_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_1 = head ? data_1_state_0_1 : data_0_state_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_2 = head ? data_1_state_0_2 : data_0_state_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_0_3 = head ? data_1_state_0_3 : data_0_state_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_0 = head ? data_1_state_1_0 : data_0_state_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_1 = head ? data_1_state_1_1 : data_0_state_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_2 = head ? data_1_state_1_2 : data_0_state_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_1_3 = head ? data_1_state_1_3 : data_0_state_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_0 = head ? data_1_state_2_0 : data_0_state_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_1 = head ? data_1_state_2_1 : data_0_state_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_2 = head ? data_1_state_2_2 : data_0_state_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_2_3 = head ? data_1_state_2_3 : data_0_state_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_0 = head ? data_1_state_3_0 : data_0_state_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_1 = head ? data_1_state_3_1 : data_0_state_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_2 = head ? data_1_state_3_2 : data_0_state_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_state_3_3 = head ? data_1_state_3_3 : data_0_state_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire [7:0] input_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  wire  _GEN_65 = tail ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:23 AES_PipelinedElasticBuffer.scala 158:23]
  wire  _GEN_206 = ~tail; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_66 = ~tail | full_0; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_67 = tail | full_1; // @[AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 159:16 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_132 = io_in_valid & ~_GEN_65 ? _GEN_66 : full_0; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_133 = io_in_valid & ~_GEN_65 ? _GEN_67 : full_1; // @[AES_PipelinedElasticBuffer.scala 158:36 AES_PipelinedElasticBuffer.scala 150:21]
  wire  _GEN_200 = head ? full_1 : full_0; // @[AES_PipelinedElasticBuffer.scala 165:21 AES_PipelinedElasticBuffer.scala 165:21]
  AES_SubBytes sub ( // @[AES_PipelinedElasticBuffer.scala 171:19]
    .io_out_state_0_0(sub_io_out_state_0_0),
    .io_out_state_0_1(sub_io_out_state_0_1),
    .io_out_state_0_2(sub_io_out_state_0_2),
    .io_out_state_0_3(sub_io_out_state_0_3),
    .io_out_state_1_0(sub_io_out_state_1_0),
    .io_out_state_1_1(sub_io_out_state_1_1),
    .io_out_state_1_2(sub_io_out_state_1_2),
    .io_out_state_1_3(sub_io_out_state_1_3),
    .io_out_state_2_0(sub_io_out_state_2_0),
    .io_out_state_2_1(sub_io_out_state_2_1),
    .io_out_state_2_2(sub_io_out_state_2_2),
    .io_out_state_2_3(sub_io_out_state_2_3),
    .io_out_state_3_0(sub_io_out_state_3_0),
    .io_out_state_3_1(sub_io_out_state_3_1),
    .io_out_state_3_2(sub_io_out_state_3_2),
    .io_out_state_3_3(sub_io_out_state_3_3),
    .io_in_state_0_0(sub_io_in_state_0_0),
    .io_in_state_0_1(sub_io_in_state_0_1),
    .io_in_state_0_2(sub_io_in_state_0_2),
    .io_in_state_0_3(sub_io_in_state_0_3),
    .io_in_state_1_0(sub_io_in_state_1_0),
    .io_in_state_1_1(sub_io_in_state_1_1),
    .io_in_state_1_2(sub_io_in_state_1_2),
    .io_in_state_1_3(sub_io_in_state_1_3),
    .io_in_state_2_0(sub_io_in_state_2_0),
    .io_in_state_2_1(sub_io_in_state_2_1),
    .io_in_state_2_2(sub_io_in_state_2_2),
    .io_in_state_2_3(sub_io_in_state_2_3),
    .io_in_state_3_0(sub_io_in_state_3_0),
    .io_in_state_3_1(sub_io_in_state_3_1),
    .io_in_state_3_2(sub_io_in_state_3_2),
    .io_in_state_3_3(sub_io_in_state_3_3)
  );
  AES_ShiftRows shift ( // @[AES_PipelinedElasticBuffer.scala 179:21]
    .io_out_state_0_0(shift_io_out_state_0_0),
    .io_out_state_0_1(shift_io_out_state_0_1),
    .io_out_state_0_2(shift_io_out_state_0_2),
    .io_out_state_0_3(shift_io_out_state_0_3),
    .io_out_state_1_0(shift_io_out_state_1_0),
    .io_out_state_1_1(shift_io_out_state_1_1),
    .io_out_state_1_2(shift_io_out_state_1_2),
    .io_out_state_1_3(shift_io_out_state_1_3),
    .io_out_state_2_0(shift_io_out_state_2_0),
    .io_out_state_2_1(shift_io_out_state_2_1),
    .io_out_state_2_2(shift_io_out_state_2_2),
    .io_out_state_2_3(shift_io_out_state_2_3),
    .io_out_state_3_0(shift_io_out_state_3_0),
    .io_out_state_3_1(shift_io_out_state_3_1),
    .io_out_state_3_2(shift_io_out_state_3_2),
    .io_out_state_3_3(shift_io_out_state_3_3),
    .io_in_state_0_0(shift_io_in_state_0_0),
    .io_in_state_0_1(shift_io_in_state_0_1),
    .io_in_state_0_2(shift_io_in_state_0_2),
    .io_in_state_0_3(shift_io_in_state_0_3),
    .io_in_state_1_0(shift_io_in_state_1_0),
    .io_in_state_1_1(shift_io_in_state_1_1),
    .io_in_state_1_2(shift_io_in_state_1_2),
    .io_in_state_1_3(shift_io_in_state_1_3),
    .io_in_state_2_0(shift_io_in_state_2_0),
    .io_in_state_2_1(shift_io_in_state_2_1),
    .io_in_state_2_2(shift_io_in_state_2_2),
    .io_in_state_2_3(shift_io_in_state_2_3),
    .io_in_state_3_0(shift_io_in_state_3_0),
    .io_in_state_3_1(shift_io_in_state_3_1),
    .io_in_state_3_2(shift_io_in_state_3_2),
    .io_in_state_3_3(shift_io_in_state_3_3)
  );
  AES_MixColumns mix ( // @[AES_PipelinedElasticBuffer.scala 182:19]
    .io_out_state_0_0(mix_io_out_state_0_0),
    .io_out_state_0_1(mix_io_out_state_0_1),
    .io_out_state_0_2(mix_io_out_state_0_2),
    .io_out_state_0_3(mix_io_out_state_0_3),
    .io_out_state_1_0(mix_io_out_state_1_0),
    .io_out_state_1_1(mix_io_out_state_1_1),
    .io_out_state_1_2(mix_io_out_state_1_2),
    .io_out_state_1_3(mix_io_out_state_1_3),
    .io_out_state_2_0(mix_io_out_state_2_0),
    .io_out_state_2_1(mix_io_out_state_2_1),
    .io_out_state_2_2(mix_io_out_state_2_2),
    .io_out_state_2_3(mix_io_out_state_2_3),
    .io_out_state_3_0(mix_io_out_state_3_0),
    .io_out_state_3_1(mix_io_out_state_3_1),
    .io_out_state_3_2(mix_io_out_state_3_2),
    .io_out_state_3_3(mix_io_out_state_3_3),
    .io_in_state_0_0(mix_io_in_state_0_0),
    .io_in_state_0_1(mix_io_in_state_0_1),
    .io_in_state_0_2(mix_io_in_state_0_2),
    .io_in_state_0_3(mix_io_in_state_0_3),
    .io_in_state_1_0(mix_io_in_state_1_0),
    .io_in_state_1_1(mix_io_in_state_1_1),
    .io_in_state_1_2(mix_io_in_state_1_2),
    .io_in_state_1_3(mix_io_in_state_1_3),
    .io_in_state_2_0(mix_io_in_state_2_0),
    .io_in_state_2_1(mix_io_in_state_2_1),
    .io_in_state_2_2(mix_io_in_state_2_2),
    .io_in_state_2_3(mix_io_in_state_2_3),
    .io_in_state_3_0(mix_io_in_state_3_0),
    .io_in_state_3_1(mix_io_in_state_3_1),
    .io_in_state_3_2(mix_io_in_state_3_2),
    .io_in_state_3_3(mix_io_in_state_3_3)
  );
  AES_GetNewKey_9 key ( // @[AES_PipelinedElasticBuffer.scala 191:19]
    .io_out_key_0_0(key_io_out_key_0_0),
    .io_out_key_0_1(key_io_out_key_0_1),
    .io_out_key_0_2(key_io_out_key_0_2),
    .io_out_key_0_3(key_io_out_key_0_3),
    .io_out_key_1_0(key_io_out_key_1_0),
    .io_out_key_1_1(key_io_out_key_1_1),
    .io_out_key_1_2(key_io_out_key_1_2),
    .io_out_key_1_3(key_io_out_key_1_3),
    .io_out_key_2_0(key_io_out_key_2_0),
    .io_out_key_2_1(key_io_out_key_2_1),
    .io_out_key_2_2(key_io_out_key_2_2),
    .io_out_key_2_3(key_io_out_key_2_3),
    .io_out_key_3_0(key_io_out_key_3_0),
    .io_out_key_3_1(key_io_out_key_3_1),
    .io_out_key_3_2(key_io_out_key_3_2),
    .io_out_key_3_3(key_io_out_key_3_3),
    .io_in_key_0_0(key_io_in_key_0_0),
    .io_in_key_0_1(key_io_in_key_0_1),
    .io_in_key_0_2(key_io_in_key_0_2),
    .io_in_key_0_3(key_io_in_key_0_3),
    .io_in_key_1_0(key_io_in_key_1_0),
    .io_in_key_1_1(key_io_in_key_1_1),
    .io_in_key_1_2(key_io_in_key_1_2),
    .io_in_key_1_3(key_io_in_key_1_3),
    .io_in_key_2_0(key_io_in_key_2_0),
    .io_in_key_2_1(key_io_in_key_2_1),
    .io_in_key_2_2(key_io_in_key_2_2),
    .io_in_key_2_3(key_io_in_key_2_3),
    .io_in_key_3_0(key_io_in_key_3_0),
    .io_in_key_3_1(key_io_in_key_3_1),
    .io_in_key_3_2(key_io_in_key_3_2),
    .io_in_key_3_3(key_io_in_key_3_3)
  );
  assign io_out_valid = full_0 | full_1; // @[AES_PipelinedElasticBuffer.scala 153:27]
  assign io_out_bits_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_0 = key_io_out_key_0_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_1 = key_io_out_key_0_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_2 = key_io_out_key_0_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_0_3 = key_io_out_key_0_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_0 = key_io_out_key_1_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_1 = key_io_out_key_1_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_2 = key_io_out_key_1_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_1_3 = key_io_out_key_1_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_0 = key_io_out_key_2_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_1 = key_io_out_key_2_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_2 = key_io_out_key_2_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_2_3 = key_io_out_key_2_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_0 = key_io_out_key_3_0; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_1 = key_io_out_key_3_1; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_2 = key_io_out_key_3_2; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_out_bits_key_3_3 = key_io_out_key_3_3; // @[AES_PipelinedElasticBuffer.scala 154:15]
  assign io_in_ready = ~(full_0 & full_1); // @[AES_PipelinedElasticBuffer.scala 152:18]
  assign sub_io_in_state_0_0 = input_state_0_0 ^ input_key_0_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_1 = input_state_0_1 ^ input_key_0_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_2 = input_state_0_2 ^ input_key_0_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_0_3 = input_state_0_3 ^ input_key_0_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_0 = input_state_1_0 ^ input_key_1_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_1 = input_state_1_1 ^ input_key_1_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_2 = input_state_1_2 ^ input_key_1_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_1_3 = input_state_1_3 ^ input_key_1_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_0 = input_state_2_0 ^ input_key_2_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_1 = input_state_2_1 ^ input_key_2_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_2 = input_state_2_2 ^ input_key_2_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_2_3 = input_state_2_3 ^ input_key_2_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_0 = input_state_3_0 ^ input_key_3_0; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_1 = input_state_3_1 ^ input_key_3_1; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_2 = input_state_3_2 ^ input_key_3_2; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign sub_io_in_state_3_3 = input_state_3_3 ^ input_key_3_3; // @[AES_PipelinedElasticBuffer.scala 175:50]
  assign shift_io_in_state_0_0 = sub_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_1 = sub_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_2 = sub_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_0_3 = sub_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_0 = sub_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_1 = sub_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_2 = sub_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_1_3 = sub_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_0 = sub_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_1 = sub_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_2 = sub_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_2_3 = sub_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_0 = sub_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_1 = sub_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_2 = sub_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign shift_io_in_state_3_3 = sub_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 180:15]
  assign mix_io_in_state_0_0 = shift_io_out_state_0_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_1 = shift_io_out_state_0_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_2 = shift_io_out_state_0_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_0_3 = shift_io_out_state_0_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_0 = shift_io_out_state_1_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_1 = shift_io_out_state_1_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_2 = shift_io_out_state_1_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_1_3 = shift_io_out_state_1_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_0 = shift_io_out_state_2_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_1 = shift_io_out_state_2_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_2 = shift_io_out_state_2_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_2_3 = shift_io_out_state_2_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_0 = shift_io_out_state_3_0; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_1 = shift_io_out_state_3_1; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_2 = shift_io_out_state_3_2; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign mix_io_in_state_3_3 = shift_io_out_state_3_3; // @[AES_PipelinedElasticBuffer.scala 183:13]
  assign key_io_in_key_0_0 = head ? data_1_key_0_0 : data_0_key_0_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_1 = head ? data_1_key_0_1 : data_0_key_0_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_2 = head ? data_1_key_0_2 : data_0_key_0_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_0_3 = head ? data_1_key_0_3 : data_0_key_0_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_0 = head ? data_1_key_1_0 : data_0_key_1_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_1 = head ? data_1_key_1_1 : data_0_key_1_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_2 = head ? data_1_key_1_2 : data_0_key_1_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_1_3 = head ? data_1_key_1_3 : data_0_key_1_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_0 = head ? data_1_key_2_0 : data_0_key_2_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_1 = head ? data_1_key_2_1 : data_0_key_2_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_2 = head ? data_1_key_2_2 : data_0_key_2_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_2_3 = head ? data_1_key_2_3 : data_0_key_2_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_0 = head ? data_1_key_3_0 : data_0_key_3_0; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_1 = head ? data_1_key_3_1 : data_0_key_3_1; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_2 = head ? data_1_key_3_2 : data_0_key_3_2; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  assign key_io_in_key_3_3 = head ? data_1_key_3_3 : data_0_key_3_3; // @[AES_PipelinedElasticBuffer.scala 155:9 AES_PipelinedElasticBuffer.scala 155:9]
  always @(posedge clock) begin
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_0_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (~tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_0_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_0 <= io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_1 <= io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_2 <= io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_0_3 <= io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_0 <= io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_1 <= io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_2 <= io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_1_3 <= io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_0 <= io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_1 <= io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_2 <= io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_2_3 <= io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_0 <= io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_1 <= io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_2 <= io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_state_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_state_3_3 <= io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_0 <= io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_1 <= io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_2 <= io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_0_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_0_3 <= io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_0 <= io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_1 <= io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_2 <= io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_1_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_1_3 <= io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_0 <= io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_1 <= io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_2 <= io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_2_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_2_3 <= io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_0 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_0 <= io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_1 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_1 <= io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_2 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_2 <= io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 147:21]
      data_1_key_3_3 <= 8'h0; // @[AES_PipelinedElasticBuffer.scala 147:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      if (tail) begin // @[AES_PipelinedElasticBuffer.scala 160:16]
        data_1_key_3_3 <= io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 160:16]
      end
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 148:21]
      head <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 148:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      head <= ~head; // @[AES_PipelinedElasticBuffer.scala 167:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 149:21]
      tail <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 149:21]
    end else if (io_in_valid & ~_GEN_65) begin // @[AES_PipelinedElasticBuffer.scala 158:36]
      tail <= _GEN_206; // @[AES_PipelinedElasticBuffer.scala 161:10]
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (~head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_0 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_0 <= _GEN_132;
      end
    end else begin
      full_0 <= _GEN_132;
    end
    if (reset) begin // @[AES_PipelinedElasticBuffer.scala 150:21]
      full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 150:21]
    end else if (io_out_ready & _GEN_200) begin // @[AES_PipelinedElasticBuffer.scala 165:36]
      if (head) begin // @[AES_PipelinedElasticBuffer.scala 166:16]
        full_1 <= 1'h0; // @[AES_PipelinedElasticBuffer.scala 166:16]
      end else begin
        full_1 <= _GEN_133;
      end
    end else begin
      full_1 <= _GEN_133;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_state_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_state_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_0_state_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_0_state_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_0_state_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_0_state_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_0_state_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_0_state_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_0_state_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_0_state_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_0_state_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_0_state_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_0_state_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_0_state_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_0_state_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_0_state_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_0_key_0_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_0_key_0_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_0_key_0_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_0_key_0_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_0_key_1_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_0_key_1_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_0_key_1_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_0_key_1_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_0_key_2_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_0_key_2_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_0_key_2_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_0_key_2_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_0_key_3_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_0_key_3_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_0_key_3_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_0_key_3_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_1_state_0_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_1_state_0_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_1_state_0_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_1_state_0_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_1_state_1_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_1_state_1_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_1_state_1_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_1_state_1_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_1_state_2_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_1_state_2_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_1_state_2_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  data_1_state_2_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  data_1_state_3_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  data_1_state_3_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  data_1_state_3_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  data_1_state_3_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  data_1_key_0_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  data_1_key_0_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  data_1_key_0_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  data_1_key_0_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  data_1_key_1_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  data_1_key_1_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  data_1_key_1_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  data_1_key_1_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  data_1_key_2_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  data_1_key_2_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  data_1_key_2_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  data_1_key_2_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  data_1_key_3_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  data_1_key_3_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  data_1_key_3_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  data_1_key_3_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  head = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tail = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  full_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  full_1 = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AES_PipelinedElasticBuffer(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [127:0] io_in_bits_text,
  input  [127:0] io_in_bits_key,
  input          io_result_ready,
  output         io_result_valid,
  output [127:0] io_result_bits
);
  wire  initialPermutation_clock; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire  initialPermutation_reset; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire  initialPermutation_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire  initialPermutation_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [127:0] initialPermutation_io_in_bits_text; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [127:0] initialPermutation_io_in_bits_key; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire  initialPermutation_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire  initialPermutation_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire [7:0] initialPermutation_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 15:34]
  wire  finalPermutation_clock; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire  finalPermutation_reset; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire  finalPermutation_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire  finalPermutation_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [127:0] finalPermutation_io_out_bits; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire  finalPermutation_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire  finalPermutation_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire [7:0] finalPermutation_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 21:32]
  wire  PEs_0_clock; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_0_reset; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_0_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_0_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_0_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_0_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_0_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_1_clock; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_1_reset; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_1_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_1_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_1_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_1_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_1_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_2_clock; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_2_reset; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_2_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_2_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_2_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_2_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_2_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_3_clock; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_3_reset; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_3_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_3_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_3_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_3_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_3_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_4_clock; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_4_reset; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_4_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_4_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_4_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_4_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_4_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_5_clock; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_5_reset; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_5_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_5_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_5_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_5_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_5_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_6_clock; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_6_reset; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_6_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_6_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_6_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_6_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_6_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_7_clock; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_7_reset; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_7_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_7_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_7_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_7_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_7_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_8_clock; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_8_reset; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_8_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_8_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_8_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_8_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_8_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_9_clock; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_9_reset; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_9_io_out_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_9_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_9_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire  PEs_9_io_in_valid; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 27:20]
  wire [7:0] PEs_9_io_in_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 27:20]
  AES_InitialOperation initialPermutation ( // @[AES_PipelinedElasticBuffer.scala 15:34]
    .clock(initialPermutation_clock),
    .reset(initialPermutation_reset),
    .io_in_ready(initialPermutation_io_in_ready),
    .io_in_valid(initialPermutation_io_in_valid),
    .io_in_bits_text(initialPermutation_io_in_bits_text),
    .io_in_bits_key(initialPermutation_io_in_bits_key),
    .io_out_ready(initialPermutation_io_out_ready),
    .io_out_valid(initialPermutation_io_out_valid),
    .io_out_bits_state_0_0(initialPermutation_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(initialPermutation_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(initialPermutation_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(initialPermutation_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(initialPermutation_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(initialPermutation_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(initialPermutation_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(initialPermutation_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(initialPermutation_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(initialPermutation_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(initialPermutation_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(initialPermutation_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(initialPermutation_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(initialPermutation_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(initialPermutation_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(initialPermutation_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(initialPermutation_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(initialPermutation_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(initialPermutation_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(initialPermutation_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(initialPermutation_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(initialPermutation_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(initialPermutation_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(initialPermutation_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(initialPermutation_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(initialPermutation_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(initialPermutation_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(initialPermutation_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(initialPermutation_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(initialPermutation_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(initialPermutation_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(initialPermutation_io_out_bits_key_3_3)
  );
  AES_FinalOperation finalPermutation ( // @[AES_PipelinedElasticBuffer.scala 21:32]
    .clock(finalPermutation_clock),
    .reset(finalPermutation_reset),
    .io_out_ready(finalPermutation_io_out_ready),
    .io_out_valid(finalPermutation_io_out_valid),
    .io_out_bits(finalPermutation_io_out_bits),
    .io_in_ready(finalPermutation_io_in_ready),
    .io_in_valid(finalPermutation_io_in_valid),
    .io_in_bits_state_0_0(finalPermutation_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(finalPermutation_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(finalPermutation_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(finalPermutation_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(finalPermutation_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(finalPermutation_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(finalPermutation_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(finalPermutation_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(finalPermutation_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(finalPermutation_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(finalPermutation_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(finalPermutation_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(finalPermutation_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(finalPermutation_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(finalPermutation_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(finalPermutation_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(finalPermutation_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(finalPermutation_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(finalPermutation_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(finalPermutation_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(finalPermutation_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(finalPermutation_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(finalPermutation_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(finalPermutation_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(finalPermutation_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(finalPermutation_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(finalPermutation_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(finalPermutation_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(finalPermutation_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(finalPermutation_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(finalPermutation_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(finalPermutation_io_in_bits_key_3_3)
  );
  AES_ProcessingElement PEs_0 ( // @[AES_PipelinedElasticBuffer.scala 27:20]
    .clock(PEs_0_clock),
    .reset(PEs_0_reset),
    .io_out_ready(PEs_0_io_out_ready),
    .io_out_valid(PEs_0_io_out_valid),
    .io_out_bits_state_0_0(PEs_0_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_0_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_0_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_0_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_0_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_0_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_0_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_0_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_0_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_0_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_0_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_0_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_0_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_0_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_0_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_0_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_0_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_0_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_0_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_0_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_0_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_0_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_0_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_0_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_0_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_0_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_0_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_0_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_0_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_0_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_0_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_0_io_out_bits_key_3_3),
    .io_in_ready(PEs_0_io_in_ready),
    .io_in_valid(PEs_0_io_in_valid),
    .io_in_bits_state_0_0(PEs_0_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_0_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_0_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_0_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_0_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_0_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_0_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_0_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_0_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_0_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_0_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_0_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_0_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_0_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_0_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_0_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_0_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_0_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_0_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_0_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_0_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_0_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_0_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_0_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_0_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_0_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_0_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_0_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_0_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_0_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_0_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_0_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_1 PEs_1 ( // @[AES_PipelinedElasticBuffer.scala 27:20]
    .clock(PEs_1_clock),
    .reset(PEs_1_reset),
    .io_out_ready(PEs_1_io_out_ready),
    .io_out_valid(PEs_1_io_out_valid),
    .io_out_bits_state_0_0(PEs_1_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_1_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_1_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_1_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_1_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_1_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_1_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_1_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_1_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_1_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_1_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_1_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_1_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_1_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_1_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_1_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_1_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_1_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_1_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_1_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_1_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_1_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_1_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_1_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_1_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_1_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_1_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_1_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_1_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_1_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_1_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_1_io_out_bits_key_3_3),
    .io_in_ready(PEs_1_io_in_ready),
    .io_in_valid(PEs_1_io_in_valid),
    .io_in_bits_state_0_0(PEs_1_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_1_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_1_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_1_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_1_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_1_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_1_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_1_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_1_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_1_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_1_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_1_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_1_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_1_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_1_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_1_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_1_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_1_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_1_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_1_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_1_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_1_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_1_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_1_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_1_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_1_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_1_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_1_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_1_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_1_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_1_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_1_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_2 PEs_2 ( // @[AES_PipelinedElasticBuffer.scala 27:20]
    .clock(PEs_2_clock),
    .reset(PEs_2_reset),
    .io_out_ready(PEs_2_io_out_ready),
    .io_out_valid(PEs_2_io_out_valid),
    .io_out_bits_state_0_0(PEs_2_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_2_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_2_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_2_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_2_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_2_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_2_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_2_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_2_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_2_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_2_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_2_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_2_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_2_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_2_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_2_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_2_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_2_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_2_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_2_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_2_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_2_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_2_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_2_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_2_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_2_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_2_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_2_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_2_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_2_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_2_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_2_io_out_bits_key_3_3),
    .io_in_ready(PEs_2_io_in_ready),
    .io_in_valid(PEs_2_io_in_valid),
    .io_in_bits_state_0_0(PEs_2_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_2_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_2_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_2_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_2_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_2_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_2_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_2_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_2_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_2_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_2_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_2_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_2_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_2_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_2_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_2_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_2_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_2_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_2_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_2_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_2_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_2_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_2_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_2_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_2_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_2_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_2_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_2_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_2_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_2_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_2_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_2_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_3 PEs_3 ( // @[AES_PipelinedElasticBuffer.scala 27:20]
    .clock(PEs_3_clock),
    .reset(PEs_3_reset),
    .io_out_ready(PEs_3_io_out_ready),
    .io_out_valid(PEs_3_io_out_valid),
    .io_out_bits_state_0_0(PEs_3_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_3_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_3_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_3_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_3_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_3_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_3_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_3_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_3_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_3_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_3_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_3_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_3_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_3_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_3_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_3_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_3_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_3_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_3_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_3_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_3_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_3_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_3_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_3_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_3_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_3_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_3_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_3_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_3_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_3_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_3_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_3_io_out_bits_key_3_3),
    .io_in_ready(PEs_3_io_in_ready),
    .io_in_valid(PEs_3_io_in_valid),
    .io_in_bits_state_0_0(PEs_3_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_3_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_3_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_3_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_3_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_3_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_3_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_3_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_3_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_3_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_3_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_3_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_3_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_3_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_3_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_3_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_3_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_3_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_3_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_3_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_3_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_3_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_3_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_3_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_3_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_3_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_3_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_3_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_3_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_3_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_3_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_3_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_4 PEs_4 ( // @[AES_PipelinedElasticBuffer.scala 27:20]
    .clock(PEs_4_clock),
    .reset(PEs_4_reset),
    .io_out_ready(PEs_4_io_out_ready),
    .io_out_valid(PEs_4_io_out_valid),
    .io_out_bits_state_0_0(PEs_4_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_4_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_4_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_4_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_4_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_4_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_4_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_4_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_4_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_4_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_4_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_4_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_4_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_4_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_4_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_4_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_4_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_4_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_4_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_4_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_4_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_4_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_4_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_4_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_4_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_4_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_4_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_4_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_4_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_4_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_4_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_4_io_out_bits_key_3_3),
    .io_in_ready(PEs_4_io_in_ready),
    .io_in_valid(PEs_4_io_in_valid),
    .io_in_bits_state_0_0(PEs_4_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_4_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_4_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_4_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_4_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_4_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_4_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_4_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_4_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_4_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_4_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_4_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_4_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_4_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_4_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_4_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_4_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_4_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_4_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_4_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_4_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_4_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_4_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_4_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_4_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_4_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_4_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_4_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_4_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_4_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_4_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_4_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_5 PEs_5 ( // @[AES_PipelinedElasticBuffer.scala 27:20]
    .clock(PEs_5_clock),
    .reset(PEs_5_reset),
    .io_out_ready(PEs_5_io_out_ready),
    .io_out_valid(PEs_5_io_out_valid),
    .io_out_bits_state_0_0(PEs_5_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_5_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_5_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_5_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_5_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_5_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_5_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_5_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_5_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_5_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_5_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_5_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_5_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_5_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_5_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_5_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_5_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_5_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_5_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_5_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_5_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_5_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_5_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_5_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_5_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_5_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_5_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_5_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_5_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_5_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_5_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_5_io_out_bits_key_3_3),
    .io_in_ready(PEs_5_io_in_ready),
    .io_in_valid(PEs_5_io_in_valid),
    .io_in_bits_state_0_0(PEs_5_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_5_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_5_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_5_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_5_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_5_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_5_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_5_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_5_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_5_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_5_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_5_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_5_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_5_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_5_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_5_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_5_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_5_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_5_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_5_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_5_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_5_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_5_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_5_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_5_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_5_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_5_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_5_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_5_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_5_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_5_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_5_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_6 PEs_6 ( // @[AES_PipelinedElasticBuffer.scala 27:20]
    .clock(PEs_6_clock),
    .reset(PEs_6_reset),
    .io_out_ready(PEs_6_io_out_ready),
    .io_out_valid(PEs_6_io_out_valid),
    .io_out_bits_state_0_0(PEs_6_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_6_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_6_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_6_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_6_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_6_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_6_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_6_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_6_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_6_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_6_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_6_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_6_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_6_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_6_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_6_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_6_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_6_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_6_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_6_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_6_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_6_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_6_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_6_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_6_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_6_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_6_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_6_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_6_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_6_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_6_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_6_io_out_bits_key_3_3),
    .io_in_ready(PEs_6_io_in_ready),
    .io_in_valid(PEs_6_io_in_valid),
    .io_in_bits_state_0_0(PEs_6_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_6_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_6_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_6_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_6_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_6_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_6_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_6_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_6_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_6_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_6_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_6_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_6_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_6_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_6_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_6_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_6_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_6_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_6_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_6_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_6_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_6_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_6_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_6_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_6_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_6_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_6_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_6_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_6_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_6_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_6_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_6_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_7 PEs_7 ( // @[AES_PipelinedElasticBuffer.scala 27:20]
    .clock(PEs_7_clock),
    .reset(PEs_7_reset),
    .io_out_ready(PEs_7_io_out_ready),
    .io_out_valid(PEs_7_io_out_valid),
    .io_out_bits_state_0_0(PEs_7_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_7_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_7_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_7_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_7_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_7_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_7_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_7_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_7_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_7_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_7_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_7_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_7_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_7_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_7_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_7_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_7_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_7_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_7_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_7_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_7_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_7_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_7_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_7_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_7_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_7_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_7_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_7_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_7_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_7_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_7_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_7_io_out_bits_key_3_3),
    .io_in_ready(PEs_7_io_in_ready),
    .io_in_valid(PEs_7_io_in_valid),
    .io_in_bits_state_0_0(PEs_7_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_7_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_7_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_7_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_7_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_7_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_7_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_7_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_7_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_7_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_7_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_7_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_7_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_7_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_7_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_7_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_7_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_7_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_7_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_7_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_7_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_7_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_7_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_7_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_7_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_7_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_7_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_7_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_7_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_7_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_7_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_7_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_8 PEs_8 ( // @[AES_PipelinedElasticBuffer.scala 27:20]
    .clock(PEs_8_clock),
    .reset(PEs_8_reset),
    .io_out_ready(PEs_8_io_out_ready),
    .io_out_valid(PEs_8_io_out_valid),
    .io_out_bits_state_0_0(PEs_8_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_8_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_8_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_8_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_8_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_8_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_8_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_8_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_8_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_8_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_8_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_8_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_8_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_8_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_8_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_8_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_8_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_8_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_8_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_8_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_8_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_8_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_8_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_8_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_8_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_8_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_8_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_8_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_8_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_8_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_8_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_8_io_out_bits_key_3_3),
    .io_in_ready(PEs_8_io_in_ready),
    .io_in_valid(PEs_8_io_in_valid),
    .io_in_bits_state_0_0(PEs_8_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_8_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_8_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_8_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_8_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_8_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_8_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_8_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_8_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_8_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_8_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_8_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_8_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_8_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_8_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_8_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_8_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_8_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_8_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_8_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_8_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_8_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_8_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_8_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_8_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_8_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_8_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_8_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_8_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_8_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_8_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_8_io_in_bits_key_3_3)
  );
  AES_ProcessingElement_9 PEs_9 ( // @[AES_PipelinedElasticBuffer.scala 27:20]
    .clock(PEs_9_clock),
    .reset(PEs_9_reset),
    .io_out_ready(PEs_9_io_out_ready),
    .io_out_valid(PEs_9_io_out_valid),
    .io_out_bits_state_0_0(PEs_9_io_out_bits_state_0_0),
    .io_out_bits_state_0_1(PEs_9_io_out_bits_state_0_1),
    .io_out_bits_state_0_2(PEs_9_io_out_bits_state_0_2),
    .io_out_bits_state_0_3(PEs_9_io_out_bits_state_0_3),
    .io_out_bits_state_1_0(PEs_9_io_out_bits_state_1_0),
    .io_out_bits_state_1_1(PEs_9_io_out_bits_state_1_1),
    .io_out_bits_state_1_2(PEs_9_io_out_bits_state_1_2),
    .io_out_bits_state_1_3(PEs_9_io_out_bits_state_1_3),
    .io_out_bits_state_2_0(PEs_9_io_out_bits_state_2_0),
    .io_out_bits_state_2_1(PEs_9_io_out_bits_state_2_1),
    .io_out_bits_state_2_2(PEs_9_io_out_bits_state_2_2),
    .io_out_bits_state_2_3(PEs_9_io_out_bits_state_2_3),
    .io_out_bits_state_3_0(PEs_9_io_out_bits_state_3_0),
    .io_out_bits_state_3_1(PEs_9_io_out_bits_state_3_1),
    .io_out_bits_state_3_2(PEs_9_io_out_bits_state_3_2),
    .io_out_bits_state_3_3(PEs_9_io_out_bits_state_3_3),
    .io_out_bits_key_0_0(PEs_9_io_out_bits_key_0_0),
    .io_out_bits_key_0_1(PEs_9_io_out_bits_key_0_1),
    .io_out_bits_key_0_2(PEs_9_io_out_bits_key_0_2),
    .io_out_bits_key_0_3(PEs_9_io_out_bits_key_0_3),
    .io_out_bits_key_1_0(PEs_9_io_out_bits_key_1_0),
    .io_out_bits_key_1_1(PEs_9_io_out_bits_key_1_1),
    .io_out_bits_key_1_2(PEs_9_io_out_bits_key_1_2),
    .io_out_bits_key_1_3(PEs_9_io_out_bits_key_1_3),
    .io_out_bits_key_2_0(PEs_9_io_out_bits_key_2_0),
    .io_out_bits_key_2_1(PEs_9_io_out_bits_key_2_1),
    .io_out_bits_key_2_2(PEs_9_io_out_bits_key_2_2),
    .io_out_bits_key_2_3(PEs_9_io_out_bits_key_2_3),
    .io_out_bits_key_3_0(PEs_9_io_out_bits_key_3_0),
    .io_out_bits_key_3_1(PEs_9_io_out_bits_key_3_1),
    .io_out_bits_key_3_2(PEs_9_io_out_bits_key_3_2),
    .io_out_bits_key_3_3(PEs_9_io_out_bits_key_3_3),
    .io_in_ready(PEs_9_io_in_ready),
    .io_in_valid(PEs_9_io_in_valid),
    .io_in_bits_state_0_0(PEs_9_io_in_bits_state_0_0),
    .io_in_bits_state_0_1(PEs_9_io_in_bits_state_0_1),
    .io_in_bits_state_0_2(PEs_9_io_in_bits_state_0_2),
    .io_in_bits_state_0_3(PEs_9_io_in_bits_state_0_3),
    .io_in_bits_state_1_0(PEs_9_io_in_bits_state_1_0),
    .io_in_bits_state_1_1(PEs_9_io_in_bits_state_1_1),
    .io_in_bits_state_1_2(PEs_9_io_in_bits_state_1_2),
    .io_in_bits_state_1_3(PEs_9_io_in_bits_state_1_3),
    .io_in_bits_state_2_0(PEs_9_io_in_bits_state_2_0),
    .io_in_bits_state_2_1(PEs_9_io_in_bits_state_2_1),
    .io_in_bits_state_2_2(PEs_9_io_in_bits_state_2_2),
    .io_in_bits_state_2_3(PEs_9_io_in_bits_state_2_3),
    .io_in_bits_state_3_0(PEs_9_io_in_bits_state_3_0),
    .io_in_bits_state_3_1(PEs_9_io_in_bits_state_3_1),
    .io_in_bits_state_3_2(PEs_9_io_in_bits_state_3_2),
    .io_in_bits_state_3_3(PEs_9_io_in_bits_state_3_3),
    .io_in_bits_key_0_0(PEs_9_io_in_bits_key_0_0),
    .io_in_bits_key_0_1(PEs_9_io_in_bits_key_0_1),
    .io_in_bits_key_0_2(PEs_9_io_in_bits_key_0_2),
    .io_in_bits_key_0_3(PEs_9_io_in_bits_key_0_3),
    .io_in_bits_key_1_0(PEs_9_io_in_bits_key_1_0),
    .io_in_bits_key_1_1(PEs_9_io_in_bits_key_1_1),
    .io_in_bits_key_1_2(PEs_9_io_in_bits_key_1_2),
    .io_in_bits_key_1_3(PEs_9_io_in_bits_key_1_3),
    .io_in_bits_key_2_0(PEs_9_io_in_bits_key_2_0),
    .io_in_bits_key_2_1(PEs_9_io_in_bits_key_2_1),
    .io_in_bits_key_2_2(PEs_9_io_in_bits_key_2_2),
    .io_in_bits_key_2_3(PEs_9_io_in_bits_key_2_3),
    .io_in_bits_key_3_0(PEs_9_io_in_bits_key_3_0),
    .io_in_bits_key_3_1(PEs_9_io_in_bits_key_3_1),
    .io_in_bits_key_3_2(PEs_9_io_in_bits_key_3_2),
    .io_in_bits_key_3_3(PEs_9_io_in_bits_key_3_3)
  );
  assign io_in_ready = initialPermutation_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 19:15]
  assign io_result_valid = finalPermutation_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 23:19]
  assign io_result_bits = finalPermutation_io_out_bits; // @[AES_PipelinedElasticBuffer.scala 22:18]
  assign initialPermutation_clock = clock;
  assign initialPermutation_reset = reset;
  assign initialPermutation_io_in_valid = io_in_valid; // @[AES_PipelinedElasticBuffer.scala 16:34]
  assign initialPermutation_io_in_bits_text = io_in_bits_text; // @[AES_PipelinedElasticBuffer.scala 17:38]
  assign initialPermutation_io_in_bits_key = io_in_bits_key; // @[AES_PipelinedElasticBuffer.scala 18:37]
  assign initialPermutation_io_out_ready = PEs_0_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 36:39]
  assign finalPermutation_clock = clock;
  assign finalPermutation_reset = reset;
  assign finalPermutation_io_out_ready = io_result_ready; // @[AES_PipelinedElasticBuffer.scala 24:33]
  assign finalPermutation_io_in_valid = PEs_9_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 42:36]
  assign finalPermutation_io_in_bits_state_0_0 = PEs_9_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_0_1 = PEs_9_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_0_2 = PEs_9_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_0_3 = PEs_9_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_1_0 = PEs_9_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_1_1 = PEs_9_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_1_2 = PEs_9_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_1_3 = PEs_9_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_2_0 = PEs_9_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_2_1 = PEs_9_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_2_2 = PEs_9_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_2_3 = PEs_9_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_3_0 = PEs_9_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_3_1 = PEs_9_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_3_2 = PEs_9_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_state_3_3 = PEs_9_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 43:41]
  assign finalPermutation_io_in_bits_key_0_0 = PEs_9_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_0_1 = PEs_9_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_0_2 = PEs_9_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_0_3 = PEs_9_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_1_0 = PEs_9_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_1_1 = PEs_9_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_1_2 = PEs_9_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_1_3 = PEs_9_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_2_0 = PEs_9_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_2_1 = PEs_9_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_2_2 = PEs_9_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_2_3 = PEs_9_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_3_0 = PEs_9_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_3_1 = PEs_9_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_3_2 = PEs_9_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign finalPermutation_io_in_bits_key_3_3 = PEs_9_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 44:39]
  assign PEs_0_clock = clock;
  assign PEs_0_reset = reset;
  assign PEs_0_io_out_ready = PEs_1_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 40:27]
  assign PEs_0_io_in_valid = initialPermutation_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 34:26]
  assign PEs_0_io_in_bits_state_0_0 = initialPermutation_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_0_1 = initialPermutation_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_0_2 = initialPermutation_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_0_3 = initialPermutation_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_1_0 = initialPermutation_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_1_1 = initialPermutation_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_1_2 = initialPermutation_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_1_3 = initialPermutation_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_2_0 = initialPermutation_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_2_1 = initialPermutation_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_2_2 = initialPermutation_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_2_3 = initialPermutation_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_3_0 = initialPermutation_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_3_1 = initialPermutation_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_3_2 = initialPermutation_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_state_3_3 = initialPermutation_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_0_0 = initialPermutation_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_0_1 = initialPermutation_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_0_2 = initialPermutation_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_0_3 = initialPermutation_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_1_0 = initialPermutation_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_1_1 = initialPermutation_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_1_2 = initialPermutation_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_1_3 = initialPermutation_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_2_0 = initialPermutation_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_2_1 = initialPermutation_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_2_2 = initialPermutation_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_2_3 = initialPermutation_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_3_0 = initialPermutation_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_3_1 = initialPermutation_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_3_2 = initialPermutation_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_0_io_in_bits_key_3_3 = initialPermutation_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 35:25]
  assign PEs_1_clock = clock;
  assign PEs_1_reset = reset;
  assign PEs_1_io_out_ready = PEs_2_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 49:27]
  assign PEs_1_io_in_valid = PEs_0_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 38:28]
  assign PEs_1_io_in_bits_state_0_0 = PEs_0_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_0_1 = PEs_0_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_0_2 = PEs_0_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_0_3 = PEs_0_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_1_0 = PEs_0_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_1_1 = PEs_0_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_1_2 = PEs_0_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_1_3 = PEs_0_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_2_0 = PEs_0_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_2_1 = PEs_0_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_2_2 = PEs_0_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_2_3 = PEs_0_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_3_0 = PEs_0_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_3_1 = PEs_0_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_3_2 = PEs_0_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_state_3_3 = PEs_0_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_0_0 = PEs_0_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_0_1 = PEs_0_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_0_2 = PEs_0_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_0_3 = PEs_0_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_1_0 = PEs_0_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_1_1 = PEs_0_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_1_2 = PEs_0_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_1_3 = PEs_0_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_2_0 = PEs_0_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_2_1 = PEs_0_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_2_2 = PEs_0_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_2_3 = PEs_0_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_3_0 = PEs_0_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_3_1 = PEs_0_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_3_2 = PEs_0_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_1_io_in_bits_key_3_3 = PEs_0_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 39:27]
  assign PEs_2_clock = clock;
  assign PEs_2_reset = reset;
  assign PEs_2_io_out_ready = PEs_3_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 49:27]
  assign PEs_2_io_in_valid = PEs_1_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 47:28]
  assign PEs_2_io_in_bits_state_0_0 = PEs_1_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_0_1 = PEs_1_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_0_2 = PEs_1_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_0_3 = PEs_1_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_1_0 = PEs_1_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_1_1 = PEs_1_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_1_2 = PEs_1_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_1_3 = PEs_1_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_2_0 = PEs_1_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_2_1 = PEs_1_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_2_2 = PEs_1_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_2_3 = PEs_1_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_3_0 = PEs_1_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_3_1 = PEs_1_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_3_2 = PEs_1_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_state_3_3 = PEs_1_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_0_0 = PEs_1_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_0_1 = PEs_1_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_0_2 = PEs_1_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_0_3 = PEs_1_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_1_0 = PEs_1_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_1_1 = PEs_1_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_1_2 = PEs_1_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_1_3 = PEs_1_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_2_0 = PEs_1_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_2_1 = PEs_1_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_2_2 = PEs_1_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_2_3 = PEs_1_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_3_0 = PEs_1_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_3_1 = PEs_1_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_3_2 = PEs_1_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_2_io_in_bits_key_3_3 = PEs_1_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_clock = clock;
  assign PEs_3_reset = reset;
  assign PEs_3_io_out_ready = PEs_4_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 49:27]
  assign PEs_3_io_in_valid = PEs_2_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 47:28]
  assign PEs_3_io_in_bits_state_0_0 = PEs_2_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_0_1 = PEs_2_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_0_2 = PEs_2_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_0_3 = PEs_2_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_1_0 = PEs_2_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_1_1 = PEs_2_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_1_2 = PEs_2_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_1_3 = PEs_2_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_2_0 = PEs_2_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_2_1 = PEs_2_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_2_2 = PEs_2_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_2_3 = PEs_2_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_3_0 = PEs_2_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_3_1 = PEs_2_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_3_2 = PEs_2_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_state_3_3 = PEs_2_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_0_0 = PEs_2_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_0_1 = PEs_2_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_0_2 = PEs_2_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_0_3 = PEs_2_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_1_0 = PEs_2_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_1_1 = PEs_2_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_1_2 = PEs_2_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_1_3 = PEs_2_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_2_0 = PEs_2_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_2_1 = PEs_2_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_2_2 = PEs_2_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_2_3 = PEs_2_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_3_0 = PEs_2_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_3_1 = PEs_2_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_3_2 = PEs_2_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_3_io_in_bits_key_3_3 = PEs_2_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_clock = clock;
  assign PEs_4_reset = reset;
  assign PEs_4_io_out_ready = PEs_5_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 49:27]
  assign PEs_4_io_in_valid = PEs_3_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 47:28]
  assign PEs_4_io_in_bits_state_0_0 = PEs_3_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_0_1 = PEs_3_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_0_2 = PEs_3_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_0_3 = PEs_3_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_1_0 = PEs_3_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_1_1 = PEs_3_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_1_2 = PEs_3_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_1_3 = PEs_3_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_2_0 = PEs_3_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_2_1 = PEs_3_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_2_2 = PEs_3_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_2_3 = PEs_3_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_3_0 = PEs_3_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_3_1 = PEs_3_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_3_2 = PEs_3_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_state_3_3 = PEs_3_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_0_0 = PEs_3_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_0_1 = PEs_3_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_0_2 = PEs_3_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_0_3 = PEs_3_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_1_0 = PEs_3_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_1_1 = PEs_3_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_1_2 = PEs_3_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_1_3 = PEs_3_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_2_0 = PEs_3_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_2_1 = PEs_3_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_2_2 = PEs_3_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_2_3 = PEs_3_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_3_0 = PEs_3_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_3_1 = PEs_3_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_3_2 = PEs_3_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_4_io_in_bits_key_3_3 = PEs_3_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_clock = clock;
  assign PEs_5_reset = reset;
  assign PEs_5_io_out_ready = PEs_6_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 49:27]
  assign PEs_5_io_in_valid = PEs_4_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 47:28]
  assign PEs_5_io_in_bits_state_0_0 = PEs_4_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_0_1 = PEs_4_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_0_2 = PEs_4_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_0_3 = PEs_4_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_1_0 = PEs_4_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_1_1 = PEs_4_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_1_2 = PEs_4_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_1_3 = PEs_4_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_2_0 = PEs_4_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_2_1 = PEs_4_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_2_2 = PEs_4_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_2_3 = PEs_4_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_3_0 = PEs_4_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_3_1 = PEs_4_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_3_2 = PEs_4_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_state_3_3 = PEs_4_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_0_0 = PEs_4_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_0_1 = PEs_4_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_0_2 = PEs_4_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_0_3 = PEs_4_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_1_0 = PEs_4_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_1_1 = PEs_4_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_1_2 = PEs_4_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_1_3 = PEs_4_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_2_0 = PEs_4_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_2_1 = PEs_4_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_2_2 = PEs_4_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_2_3 = PEs_4_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_3_0 = PEs_4_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_3_1 = PEs_4_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_3_2 = PEs_4_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_5_io_in_bits_key_3_3 = PEs_4_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_clock = clock;
  assign PEs_6_reset = reset;
  assign PEs_6_io_out_ready = PEs_7_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 49:27]
  assign PEs_6_io_in_valid = PEs_5_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 47:28]
  assign PEs_6_io_in_bits_state_0_0 = PEs_5_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_0_1 = PEs_5_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_0_2 = PEs_5_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_0_3 = PEs_5_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_1_0 = PEs_5_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_1_1 = PEs_5_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_1_2 = PEs_5_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_1_3 = PEs_5_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_2_0 = PEs_5_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_2_1 = PEs_5_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_2_2 = PEs_5_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_2_3 = PEs_5_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_3_0 = PEs_5_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_3_1 = PEs_5_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_3_2 = PEs_5_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_state_3_3 = PEs_5_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_0_0 = PEs_5_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_0_1 = PEs_5_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_0_2 = PEs_5_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_0_3 = PEs_5_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_1_0 = PEs_5_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_1_1 = PEs_5_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_1_2 = PEs_5_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_1_3 = PEs_5_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_2_0 = PEs_5_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_2_1 = PEs_5_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_2_2 = PEs_5_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_2_3 = PEs_5_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_3_0 = PEs_5_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_3_1 = PEs_5_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_3_2 = PEs_5_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_6_io_in_bits_key_3_3 = PEs_5_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_clock = clock;
  assign PEs_7_reset = reset;
  assign PEs_7_io_out_ready = PEs_8_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 49:27]
  assign PEs_7_io_in_valid = PEs_6_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 47:28]
  assign PEs_7_io_in_bits_state_0_0 = PEs_6_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_0_1 = PEs_6_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_0_2 = PEs_6_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_0_3 = PEs_6_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_1_0 = PEs_6_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_1_1 = PEs_6_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_1_2 = PEs_6_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_1_3 = PEs_6_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_2_0 = PEs_6_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_2_1 = PEs_6_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_2_2 = PEs_6_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_2_3 = PEs_6_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_3_0 = PEs_6_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_3_1 = PEs_6_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_3_2 = PEs_6_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_state_3_3 = PEs_6_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_0_0 = PEs_6_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_0_1 = PEs_6_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_0_2 = PEs_6_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_0_3 = PEs_6_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_1_0 = PEs_6_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_1_1 = PEs_6_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_1_2 = PEs_6_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_1_3 = PEs_6_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_2_0 = PEs_6_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_2_1 = PEs_6_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_2_2 = PEs_6_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_2_3 = PEs_6_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_3_0 = PEs_6_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_3_1 = PEs_6_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_3_2 = PEs_6_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_7_io_in_bits_key_3_3 = PEs_6_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_clock = clock;
  assign PEs_8_reset = reset;
  assign PEs_8_io_out_ready = PEs_9_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 49:27]
  assign PEs_8_io_in_valid = PEs_7_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 47:28]
  assign PEs_8_io_in_bits_state_0_0 = PEs_7_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_0_1 = PEs_7_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_0_2 = PEs_7_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_0_3 = PEs_7_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_1_0 = PEs_7_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_1_1 = PEs_7_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_1_2 = PEs_7_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_1_3 = PEs_7_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_2_0 = PEs_7_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_2_1 = PEs_7_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_2_2 = PEs_7_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_2_3 = PEs_7_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_3_0 = PEs_7_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_3_1 = PEs_7_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_3_2 = PEs_7_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_state_3_3 = PEs_7_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_0_0 = PEs_7_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_0_1 = PEs_7_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_0_2 = PEs_7_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_0_3 = PEs_7_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_1_0 = PEs_7_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_1_1 = PEs_7_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_1_2 = PEs_7_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_1_3 = PEs_7_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_2_0 = PEs_7_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_2_1 = PEs_7_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_2_2 = PEs_7_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_2_3 = PEs_7_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_3_0 = PEs_7_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_3_1 = PEs_7_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_3_2 = PEs_7_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_8_io_in_bits_key_3_3 = PEs_7_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_clock = clock;
  assign PEs_9_reset = reset;
  assign PEs_9_io_out_ready = finalPermutation_io_in_ready; // @[AES_PipelinedElasticBuffer.scala 45:27]
  assign PEs_9_io_in_valid = PEs_8_io_out_valid; // @[AES_PipelinedElasticBuffer.scala 47:28]
  assign PEs_9_io_in_bits_state_0_0 = PEs_8_io_out_bits_state_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_0_1 = PEs_8_io_out_bits_state_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_0_2 = PEs_8_io_out_bits_state_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_0_3 = PEs_8_io_out_bits_state_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_1_0 = PEs_8_io_out_bits_state_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_1_1 = PEs_8_io_out_bits_state_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_1_2 = PEs_8_io_out_bits_state_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_1_3 = PEs_8_io_out_bits_state_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_2_0 = PEs_8_io_out_bits_state_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_2_1 = PEs_8_io_out_bits_state_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_2_2 = PEs_8_io_out_bits_state_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_2_3 = PEs_8_io_out_bits_state_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_3_0 = PEs_8_io_out_bits_state_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_3_1 = PEs_8_io_out_bits_state_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_3_2 = PEs_8_io_out_bits_state_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_state_3_3 = PEs_8_io_out_bits_state_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_0_0 = PEs_8_io_out_bits_key_0_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_0_1 = PEs_8_io_out_bits_key_0_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_0_2 = PEs_8_io_out_bits_key_0_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_0_3 = PEs_8_io_out_bits_key_0_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_1_0 = PEs_8_io_out_bits_key_1_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_1_1 = PEs_8_io_out_bits_key_1_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_1_2 = PEs_8_io_out_bits_key_1_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_1_3 = PEs_8_io_out_bits_key_1_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_2_0 = PEs_8_io_out_bits_key_2_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_2_1 = PEs_8_io_out_bits_key_2_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_2_2 = PEs_8_io_out_bits_key_2_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_2_3 = PEs_8_io_out_bits_key_2_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_3_0 = PEs_8_io_out_bits_key_3_0; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_3_1 = PEs_8_io_out_bits_key_3_1; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_3_2 = PEs_8_io_out_bits_key_3_2; // @[AES_PipelinedElasticBuffer.scala 48:27]
  assign PEs_9_io_in_bits_key_3_3 = PEs_8_io_out_bits_key_3_3; // @[AES_PipelinedElasticBuffer.scala 48:27]
endmodule
